BZh91AY&SY Ԋ� h߀Px��g߰����P�wm���hW6H�y0���d� �2	�I���     �MA��A�44  ��&0a0�` 2i�a"AL����2#jbd 4�f$�	E,~�m%�C!�|���"�[چZ���4���͛I������ˠ0��ݒL��6d����@m�,�����)�x�d15��S�#�;{���P�!�1���m���-:��lr�gƣ��� D�uPj��*�Q�c]"J+H!D*5���1LHB萪�sG���24�$����}f�9rY]Jo�"$U��c=؎6F@�0�����D)Г�jQ��6U�%!�2!\4Ư(��ѝ�ֺ"5��_�O52�)�N�+u+TC�]�om#�Y�*";Y�~�n��Է�ɳ[�LYT���BC���ʲ���҉7XG��a@oXMϨǌR=J$.rKc<���f�.�Y�h�	�CY���D"��r��юdHpE)[+��r�܎P�
��A4fkX�3`���d>�Yj9v�I��/3��"�{2��Ʉ	tt��|W�Db!n$���eEc̔ư�	�����b��y�bz�]�2Ze��m�Z��V���$�L��#���a�9���6��L��EӞ jw�m�(�@�S� I2p1�tL��Uf�$V!��%B�F��<���$-W-�I0�9�-�]��c��$�]�
1���*X�ԍ��f�g�+3N�(F��-
6X�4q�b�2���+ �;��"�	�l��k��c'GUV��
3�ѕ���(`���Qy�q2��P�'r.U[���f[JT$�p��������w$S�	 H� 