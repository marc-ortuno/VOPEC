BZh91AY&SYoU!I _�Px���߰����P~tF`�DI&	���jM3DF��bC@�0# #	��14�i�&�G�4  �  �`20110�L�L�=L�j�j�7��F��A�z�z���b}bJjO����	����k������V.mC�Y��p�pkN.
3���}"���(F�4���]�}e�ȕT��ւ��A�aB��+�Y���J��k_�1�8�i���*�U�#�a�H	�i#=Duѥ�2l��iz��&aH,3��^m���I,�,�ܕ���� @X $3�_��촱'��Q+hۊ�EVJ�{ 
��C��61K	�H��q�7%��0+��Ρ�s�4�e&��J�(�Z)��ڔ2�����_��=u齲h[)k>5ģb��50��U,2,�M��D��BP�y��h)��S/��ѳr����#g�i`���9�(45�}�S����m" �R���3NݎP�
���� �n�3����(Ȃ<Yk����,��dnT'���h���+�	�	zz#�=y&��\�.�ǝU#�LZ@��|eJ#������쎩Ǘ穘ln�i$��I�r�B���2	��Ǹ��\v�N��Y�F�`��nE(�aO=I������0<�5���}#-#TCU;�)�q�p�l�z	���y��X=�B��b���
��F�
����
kI�H�0�WM�iHefp욄q���F�"�I(�׷�z�4ۿ �o7�L*J�2V�eu�!��kc Zj��<r�D0�$���8��$u)K�D����3/��9t�cd�`dܗ�]��BA�T�$