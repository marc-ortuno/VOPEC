BZh91AY&SY�(�� m_�Px��g߰����   P�wwwl�i�*��&Sjb�4J{@SOPi��C&!��5L�Q��=#A�      i�55'�����Ѡ �A�4�ɓF�� �0F`$!45=�$�43S� � 3SM�bOH�@�P�&Ĥ$�-��#��F��!���7�0EcH����`TՎۢ��Ct�[%e�]�d|�r���hwsC�E�"��Q�x:�IZ� ��0@��В�K�	����}��a��>.�ڣl#e�GZ4�CLE�༨�-̛K]��|�~.#���I�W�XkyE�Q���B���@XC�2Xb�iQ0nM��FLx�Scv����9��F΢(Jd�7��ù�×�̪vd��8BH$و�n� L�:α ĵ��*��R�H�)�ɟ�:x���������~b)�<�Ȱ�ѕՔ�{�?=��,�q����dc9Y�Ff&�د����[���ҭ</y}�[�D��X�gһ�iB�#��y��g+��`�e���R���0H)�("�ƖޙtS	��L����@'�'5
أ!��f$x6��+`w�qq��?!��,��0]��� (H��)�0a�r�=i٪�v͗�d8+�	�,�*/O=c̆+�)�!|���+��Ըڤ4cL&�D�s�O0�Z�؛��)B�&V�
�>@jwKm�(�@�S�y I2p1�\L��[���e�+�j��P)�lݨC�6q�Ū���=���WHqׅ���S�ʉ�hx\���7d��!���0�N"-C��r��k��hQ��Ӫ�B�%�`��Ԫy��r,���M��#��T��!�s��*
����]aM�uE��$�O�A�_1K�fHF)��݅L˼�C7�F�K[ �^o�|���H�
�:`