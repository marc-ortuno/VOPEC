BZh91AY&SY���0 @_�Px��o߰����PX^��d�BQ3F�oMQ��F���h�� �O�$� @     ���OS#�mLF��� S�2�&d`bba0�!�&�QI���&�b�?Q��� b6�����P� �߉��%� dkq�������.��j0.�/�I�ͭ��A�pdj���q����9^6S��/Q��+WJ9A����kn�ai���H`Q#;+i!Kr	AT��A^��C��m�)�O���n�}��
.��:�,4�axy���v��� [L��<Y\�jT��\�1����\��@x�����{`y����Hp�f��ȴAqc��,��^��
*�ա
Q��V��`�Z�P����.��@�7�UTa�ִ�>��$H$�$�@��<�\G�X�JT�~*^�u�GK�dh���v�j�* �`3s*�y:a0�];�CI�	�����}~�Ӎ�	殎K/L� �z/�ˠ@#���x$m�
f�峥�x�|�ԑH�7l�9 �!4q�<��<C6��I�P�GT�jԊ��1[�H�/�_<}��q�5��B��j}o,hjg���:��V�!-k�}'.�3�rp:Gr���(@��,�D�'U��#\�ƦH��r,�G�	�M�eݍ���'n̱i`�R�ݼO}ٲ�$Ҥu�;��Ʈe]:�3����=�6���]ʷ%����mx��s)�:c�}��I�d�!��wj%{^SM�'Q��̴�J����L]�z�Z��an�� �e`�h�Ҡu��hU��d��5)1{Բ"���!;u��ToЙ(��e|��Ԍ~�),˴. ¨
wo����'���7��������C���UQ�0۬h1-V?���mxN��AmV�z�.Q\1�.aКRvgg3�DjXݎlŶ��+�D�\렝Y"}�3��ඨ��HdX��J�k ��{�J�r(*�7���)�V�