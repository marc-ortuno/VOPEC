BZh91AY&SY��T� ߀Px��w߰����P~uJ��b���M��i�A����1��L� �LL&4��)�OP�4��4Ѡ@h  �`20110�L�L�	=4�қFi�� jzM=K�'�I@���� I�~��m%�2�>3pSQ�X���0,j��i��Z�7Tg�P��"N�AŶ��V��J�5ۓ$P��=��ь�/ę}<q���!
�� �>��+�&a�5+��Ա��1�,8�����ƃ��5x�3�_�l��"��9֨
1��A'8[�Z�(���G���������s��M��kcdH��v)�2P���4�fiȘ���&C���j�{�x�6��>z����)��U��^�h<�tq�\����9x�Jg�_�w�1��������c.D��a8�S8.p-L ]��ؠ<Ɨ��H.�B�$��e�|�nB�w�W�"�D3[�UEF{������m" �R�ٸ��O��(d	}���L�ā�)���2FV�vs.&f`Í�B~���X�]A��aB^Έ��~������Io��O�c��٪���2}�l/5)Ia�+�)��#}��>+�Z;,��&�4,�w�����۰��M�0���Q�I$a9���\����Gq
n��@X�4Q�UҰ�P!L#�~�^:�Q!p�w�I���
�������5�x�hb�3��s3�U�v�rLk_��J$Y3
(G��l� ݜ�B��d��mV3�����nzaa*�Vٔ+�q+��d���ق��E���H/�B�Az��LVcE�k��k���5*f�Zsir`�[���"�(HTƪl�