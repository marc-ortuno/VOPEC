BZh91AY&SY���� iߔPx��g߰����   P�wd�:�A$�z��SƩ���@� �h %S�&��G�j4=@ �   ����=F� �4 F&��4�ɓF�� �0F`$�M���4�'�h  �LL��z��"�� ��HI����#��F���k�ꛀ�#�*���0*Տ��v�etm-q�g�!�򍢹�Ei��Hq�/��w�X�K ҊH�)"�ainAT.�T�|�"���W'��Qi�m_�w���O4�.�	����o/��.��WT�0��H�g�3�4�EF�8�I�����JչJZ�Alw��D	��셳.��#	S|� @X $3'N��o7���O**QR�7�R��Q*#$A�!A�2�2 ��2ȗIĤk� f��w�~`{�әK%W���s(�՛Y��ڵ�	�ت��A?|}��F�G��j��r#l�r]SH�Q���/)����NJ�\m{�م ��[���-�?f}K�g
��Y�i(AT�}f�T'Suh��v�3\d��)J�W��x�NL�P�%�� �X̓|BsP��2 ��Yj9��,`w�q��P�1��Y�fp�i�� (H��I�ʘ1�9m�X1�:�#�v]L�Ace�%��@� �=gqL֙�j�3cؽW�GZ�	&��GO����/����M%�$';���&R�B L)ᘀ$�8�����=�A�l�"�o(
�8�l�ti�HX�\��~�9�Ɣ�mN��r�����=�O��Y4�jG"cZw�"���Vg�g#��ۂ���ZI@�<<5��kʋ +q��d�*�Yl�QY�����1����!|jj�@L�z�s�'Aӈ�jB�"kb�3�/��	<&6�,L�b�?�-�rE8P�����