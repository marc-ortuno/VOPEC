BZh91AY&SY(��/ ~ߔPx��g߰����   P�wd���'f �E4�M�<h�S�i�z4#&���4a�0�)ꇨ=@     	L��4��    �bdɣ	�bi�L#0	
b)�i=@#M ��f�B�=� 
�K0k`}������F���k�뛀옑�ib�jjŃH���}�~�j�~�b��뫕¦��T��/$G�{���V
J�R頸�*1H(�n��3I$�*i��.Y?O]s�*	�1�W�7q*�Zy��B��ͮ3�Ԭ3*��`mfN�OCc0dsc����R�M�0��t��"A�=%G��P�s�2[��3�3�L:)f5%eN�y!		,��@��3�Gn�/К+jl�T�*l���kk�P�!�j@���4�v�V�^��cC`6�ۜ�[�k�'��O�_iO�`?_��:��=`��ߙ�H��Ub��w��Z�b8�i[�[�0����c
1r��z��=���v�s0��#����'�-j$�����a��3y�:5�p,
!���c���Yˇ`�1���D�����K�y�B]6~$Kc8��M5tQ��2�Q��\L���qy��>c�Z�f���Q4@L<ӭ�)�L	�Z��曩Wh��0���3 �p����y�b6����PHJ+f2�Z:֛d�Z`�F ��L\'&'(i���M���F��H5;��yJ$�
w� 	B(�*���ػ�k0��%����T�q@vmY5�H�f�Ո{���f{q�
�\XRK^��0��1��A�*�P�za��W�+3���Uᢶ�e��{+��	(��~J���E���M4T�d��`���C�8g�!,
���?�(�� Ϫ�?a(6�&�@��D�r�e�X���C%���PF��|�"�(HF��