BZh91AY&SY��<� _�Px��w߰����P~tF`�	%�M!�5&���4d1��s �	������`���`4��2h2 ��   s �	������`���`$HI�&M5=OP3HCA�dm5=C�t��D�(�"��A�0&�^!��n�`�4��چ�U��o�okN
3���}"�ѰL}�>Q�̕rUS�R��F3�_�2�u��z�*Xg Ax{��wġ�cL휯��i�0����d8��=T͚��3�_��$ɕ���L)('�'P�r�Tӽ�!��^�:�Z �@�t��&�vZX��D���m�b	��+����!:d�M(l��	˄U�q�7%���k�J��,�(���}�|��R��mX���X:ѡF���^x�5��`��~4ʜ�cE�*-*��X�6I��c�BP�q��i��T9�LP���kڼnB����l*C2b��}B�CQ����q]]�iR�V�ǟ3N:ܡ����O�� �)���2 ��V��r�eX#�����gW�X�]a������������Fd.D��<�>$��&LZA��ǩK	Mካ
>�>��^�5��qR4�:쩂��B���8���b�r�8��AF,�#	�0jyK�E(�aO-I�����H�!��OS=+#TCV��8vo���z����L<��*7F*��5��;w�4��9�*�;R<ɍts�f��Y3T�#��m
6Ut�H!@�6=�;���f��\nƘXJ�2U�e
���6^^��hP7۫PSh��a�H/�?�H3`�9rDS\d^���|�N�E&&K ���rE8P���<�