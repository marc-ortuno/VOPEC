BZh91AY&SY�2� �ߔPx��o߰����   P�qN�&�
�%5$��MM�ѣ@ i�2MT�	�I       	L��F��&hOM��20�&�Cѓ �`A��2`�D��@S4�i�� � G��]0H}�@@ 
J���	>۽�H�0(�_��k�}��;f U�"�/Mu��scK�#�b�1c�61iF\�!�Lf��	T;�[�A�zv��T�I*�ԒӉs)xNoв�;�t�Qrr�����L�
S�+�&W$��Tc!.\o�����X�!B��_�x�����`|1��[JP�&U*�G�˙��K��o�0�6rR���1���P]y���+�R��)J���PT*7R�c@�P
�@H�j�
����M�����[�E�BA�M����B�,p��QA`�h��B&C�-U�Q؛�]�wX#/�z��)���-&%ՖGQ��������D~5s-��}dP�&�bޛ̪�*op;�<�C"������'�*�!���� j�:u�+�����;�p>N��gѠ�\��/e`fR� oNKSt����5�8cΈ�\V�i�&�{�)��;�yv��9!@t���q�(�X�)�@���R�3R�܌��0
"���ccQ�R��M�a�J lv���6���ϕKN�Ï�B�E�G �X��+����2ɖ�Ǵ��c�8�ҨO����3��D��gN��μ#|��ٮ�u�A#fj�� B����	ʚ���E���j�xa����vb�USRI��v�,�#��t�����9����Vh(ŉ �9�O	m��aO�R �d�c�?TL�1X��q�Ȳ!�΢�
a��=Y� ��B�ȷ\@�Y�D�׊�Y�nN�q��_LͶc)���;R6&5�~���t?��kP��W^�L3�6�|� g
��f�Z%]��bGSއ%D� ���MY����yx^2�P3�]aMC�¢�a�y4.~��z�ʫ2B%}nmUΓ}�41�ƙ��`��?����"�(Hq�G��