BZh91AY&SYm�7 k_�Px��g߰����   P�wd�8"U�	$S�Ц�J���MM=@��=L �F�@J�@�F��      =D%�2i�@b��C@i��&�&	��0`��$H"�"4���4dޤ�4���1'�$!��%!'���D��Kp�C[�ɸ��"�\�C�Z���ٕѬ��>b�H���EI�l&+�2��&^3��9!okE*%�G��T���*_ Hʸ?esu*!�1�+��«|#!�0�^2
��T1*a3U��\m�u쉸�qx21DX�vr)	\�+	0�E,Y��N�1d��5�M�U��1��
F��"�D�Kd�X �̝:����]��4�Q%\R ��J%�OS�`����!8�I���&�$Q�q�6;��V|;�?:��7�S��G��u�UR��vU������i�t|���U;,|�������0�=�)h�H�R��r���;��ڄ�9Sc��H2�)�h�Ǝ�3R";ѣ�IhQ��X�
Fz�~'곖m" �R���m�FuM���%ѓ� �Zֱ�3�)���Gs-ȎݦRe��.7�	�}�߷@]��� (H��G\�\�0�\9m��\:U�g�	��0o6+/O7�2�AW��0�7�Ƹ\�5C��d"B7���rbm��f� ¸z-���t�\R�D	�<0 	&N:C鉁�z�O��8�d�lCV�
a<��=Zf#p�l�zk��s[Pp�|I�������r�:v�c>�l�D���oc�"���Vg�^�'#dk3C�YWq zp֘�>9*�9i�E	Xdʍ� �R�@�)�*�ⴴ-XCI@Ӓ�����C) ͅ�~��>%0T���ܼ'c2�(S�k%���D�����H�
���