BZh91AY&SY֭`D _�Px���߰����P~tJ٦Ek����H�H���@ h�hh�&MLL`��J��MS�SCɤ     �12dф�14�&��	14�4��h�Ě  ����OH���@��� �0&�[�C[��	��i1u5
����8�w�B���N$����ʒt�'I����q���"$Ǭ�Y\g8�$[.�XdgD��J��-��[�(j��ujU]��a�l,h�pL�3a�JEnf&��WO�Izdij�`԰�IT�Ԡ=Q$�޺��tƐ����I�{߫Ɓ��4���6���FC��~Z�T� a($1od�!���^�o0�p�|3`_�����)V���<9��W�|.�#�ZV:�v=���=�Sݺ1oƈ��+|ݸ�\=hUO*˘��&��ؠ:U�����H-ڢB����?�3�i�E�<�a2�a�6T��2Ժ�8oJ�"��iJt�楐��rvC���t��P���(�{�]���-&b`�	�v =��/&%ӹ��r`��B�Ia�d��U���*`��$A���g!�b���G����fůe8ie��0�A��so�ar����Ô2%�FI�05;��qJ!@�S�� �d�c�?|L��U3�f)D5Q��B�F4�|7�9����L<M�+�+���D<��lm�L���L��J{���jc\;4�"��xQB5MW`Q��A�) ���[�|&��o�(�:���dǐDzeD�Lbf\�a�d
��f,AM�uE��H1�r���e��)�bC�\KҺ���I��dd�`d�o�w$S�	j�@