BZh91AY&SY(�e� i_�Px��g߰����   P�wd�9�������2j{T�J0������44� �M&
eP�     4��6��@h ���bdɣ	�bi�L#0	Mi�MhڛSF���z��B��� ��%P\Ĥ$��|���6��!����@"��R���0)j��jͳ�2�v���?�o�^+�=Iр/�N���{	���~(X>іrRbl�k���c�\�ބ�/�$b\O��NOq2�i����ʩ���@]��&��4(7t�'H.���ՉS��(�3A0S��F�s<��R4u �)riUBNzŚ$�-�y8g�J����0B�!�:u�}��-�4�Q%[��R ��J%E������
�I2e�N\"n��1�]3��5�G{��S⮜��i�����g�^�G��M%�m:.��2a�`}K>�{|6g�H��}kTj�M	�圕�5(^�"ɘ�o�*��~�lPU��q}�[�D��$��o0Ըԅ�GJ3}p+	��إ��Z���d�u��U�C2wO9ҵKU�[z$8�)����i��bL�	�bl���؎NR҂����<�X���^`���@L���Gu�L��j��`��V��j�a9l߮��R��H��8W��kk��ǱveV�g�I���Fm�L2��{���PH@s�$QyA�.�-��@�O�� �e1�lP��-�A�2�D5Q�&
6��f�GA!lƶ�I��Վ���ϑ@�1A��a�H�����-.60�Ѥ2d�S(q�!舒3�)Q���Bm�"Z��L$�x�G��K0Ѯ�WM�<�b�|��l8���*��T*W:�|�POH�]I40��+�C�bA��N�Q�fj��b�*N�L��K�&(�����w$S�	��_�