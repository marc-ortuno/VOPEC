BZh91AY&SYd�^ �߀Px��o߰����P��8�j���$����#ƔS#M��2� ���2	        H�Bh���2i�  �zjh`20110�L�L�l@��j�4����#UC���@��� �`SIo����p�@�Eؼ-C�X�i5q�����  c!�2�pr8x(�����W�����rX]��(�J�d����Li�=���آ��*2������aZq�	$$N�����Ӌ�P������Ua��_�|�v� �KQ��7Fd�WF��(�KA��2��hI�}+hB�z�NjE�,�P��E�FS�u�h�b�"�B�PL�2�0b��Bؤ
�Ua��f�%�[��C�;��̂��r��*M«�l�\5d��7hd�ſ;a0M��G̢ݛd��r�d{��}�H �I�6��A���x�~R,MGy���.�K��#{� ����JƘ�MH ���I����!���f��CbI���DN߽qt���=����C:yv��7�?H Y��pj������RO0�-�����=OR�Eʘ��[����z��!�@y�����H.�
S.Fvt�њP� ��e�f,	�Q^�<NʑA�Q�����7��6�E)U�i9pb�&�0�'ї�B�b�.!���(Z�̆�Yd�Q��.(X��/4*�k�@z,��`XP$�p��0`"0!n$�raR��ꯦ	��=m�]��I�8�tb��%2�f����.����i@I0���X��e
���l��4� ������s���弥aO�$$���H~� `�S��A�H�!����
a9�vUX�8Xh\s`�3Q h�B�<ED�y���1h��75�&�ԍ��g��0B��WC^ʔ#lշ-�$�w�����1���M��rlA8�`F=�"#�30�Ġk�����	������}D��h�Te"Z��	ٗ�R|wJcd�L�\#�]��BA�W�x