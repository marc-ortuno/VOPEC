BZh91AY&SY��j6 UߔPx��o߰����   P�wd�A$�jxiM=��4ɡ���@2i���@%7�hɠ     HI6�A�@h4��  �@hɉ�	���0 �`�0�"A�?)�F#H�F#@ hi�C4�> A ��������g�"Gk�%�!�în�1�H���`U�_�s����t�����0�S���Ύ">i��Y����<��jM�
l^����,��2ܐ�*VB�p?/]o�(T4Ǹ�wo
�0�������L�1���`@�u�h�C�TtH+2�8����MeȔ�Q�9(+I�dJL�J4tw^g���ڏ.96�!		*�I �1����dkp�1!��E"�!E(h��i	0�EL� �ʄ�k1D�4q֮��)����;�j�U]���[�o��^��g�G{��<�	Z��u���螚�8̯�t�bW�n��Ij4[°����n0�3	�ĩ7[]b�)ĝ"NX4�_C(X�Ԋ�@�$ �4P2�(f(��6�vU�$Hl:R���7^�š�"��m�H'���{D�f�2k-������`d�O�l�
�y[�0��&�
9|���|bB�$��m�Bމ!~Ɂ�DJ���e���9!tb���d�����6=�ӊ�u�7�I1\ii�:yQ1p�y�Ɗ�p^T�Q�A|�5<%��H L)ݼ@L�t�퉁��K��<-�dCV�B�F�mbZ4��H[o^<Ę~�:�G]8W���1썼�2�0�T��;�8��͐�Efvm��p�]�(�p��כ�%���ݭU��^���x����L��L
+v!���BZJ���)�>�(&d@�퉲���-jb�"�"�/fZH)f�A�����(*������H�
mF�