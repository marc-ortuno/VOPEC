BZh91AY&SYN׷% i_�Px��g߰����   P�wd�8(.l$� �LԌ�SG�h �i� JL��=OQ��      ��SI��h42 � @i��&�&	��0`��$HI�F!4��=LOD� f��m�����*��%!'ۓ�D��Kx�C[�ɸق1"�.f��SU�{�.�B�#; �C�&/�N�e1bh��#�c�~>�߉��Ǒ��911dƺe�nЕ��HIR��E����UwYB�i�eOǿR��E�D��xZ��s��t�����.�2��-Jp8sR+Rv�rh>�\�����!T�ReB��qo>��tmtє�Lf�B�'�t�!� ��k��(�p��'E5)�ms\�U�]qZ�,�H�DRZ"*P��*@�l�4�#�� ��|7p��x쯉Yk2}���P�i��D����Ȫ��B������U��X�mJ�TQ����58���j�I��I[֜�*�`�`):�nR�P��3i_��P��Fo�r��s�7֨15j^�3��źm" �R�ʴ�/�S^g(dD�V~$��"1M5�(Ȃ9�]�߰�L���!���>C��Y�W�.��� (H��G\�0b"��9�eqt,O ,�4�z����Ġ4�-�����0�0l|K�z�uUN	&��GNӐL\f���Xk�F��W�FI��jwK]�(�@�S� �d�c�>�� �W���,�\CX�r��L#V�!N}9	VE��I��ђ���ѕ@�[b�?F��u�f�XRd����PG	������	:�
��c:��@�-�+��*a�.BL���#�)�B	,��FD��a<X��G��!�� �������S�����j}�e�R���c;%���L_�����w$S�	�{rP