BZh91AY&SY�H� i߀Px��g߰����P�t�c��$�S�mQ���=M� ��4h�(S�b)���44�    ��B(� 4� 4�C��L`�a4� d�@�D����h�4ЦOO)4�i���>� ��%� �'���|�i/!���t���"�^C�X��:�L����?���8J�i�D�N ��}��dg���2��#qm�Z?L�P�^�b̤��*g H�=��a��;1�?�{��U�i�aXTQ*7�Ew޲ʨ���Q��X�l���¡�bJD4�`��MG$��㒣��15T$R%X��J�G}��c��ن�V�Й���b , ��_7-nwe�Ҟj$�K��D��)D��P�S*�:��e$�l�	�(�8���Ȓ�3;�~����֫�R�:�O=2�gmԯ*t��kU�r�Ep-e��v�Ӹ�xh�`"��F�Z���w�(��4'$��T����b�]`.JS.,��u^C5B�#捿ޅ�D3)fx��*��C���z��"�+eu;r���P�
����LV3�`��N��4(�7
��&�~�+\^�>ُ�W��f���2aB_o4{g�����]ėVK&�FC̕N�!������O:��!X`�&��h��sl}k璴u�7�0�ѡ�}��L\��peEi�/*n(ő$_9�Oqĥ�
y�@L�t��D���d����H�j�2��L#���C߷A�B�z�3���ٻ���Nz��3h��wu�&��H�Lkw-�2IHefuu�B8MYhQ��AӁ ������U���dn5ԕeS��A<fmKB�F8�Ӥ�x����0o=#��8��EPj�k���A�}�$KED�PT
fK�]��B@2M#�