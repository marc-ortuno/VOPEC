BZh91AY&SY�	� ߀Px��w߰����P~t��:dV�I(�j�I�4���4 ��@��#SM0M�hi�L 24 J��@P�zF��i�   9�L�����a0CLM0$ �2�=����� ��CLS�$�A@Eb I��i.ѐ�i�7�`�EL[چMX�s��6B͵���<.�}�L�S�0���j�^���T���1m�Z1�&L�˯����HB�ER���>�c��U�"ғ�XZ]��p/�ȩ��I�Ț�X�	�j+,�P�fSEeVfr����=u���!		*�I�g���S0�#��[�7u�d�Z�&�W"	�1���L�k�P��\�6�%e-�}���}a++'���:H��S8�/"mᑰ �欵�Y�Y��i�P1��LkW6��=iO���79�.�W���R�`��r�A����Is����wԅ�ތ�y��f�)f9X��/?͞��P��4�:g��l#�};!�C�S��+�3h���d>��s����?Ë�*��M�ac���}�RaB^N����F-�kK��O���T�� �Dm�l(�22ъk	��*q��5�V$ᥖK#L �P9w�0����Ӡ1�
1`I�<��.��Q
�HI������0/W�T��+�TCU
)�lߨCї1�$-���D�w�1��
�W�QA+��;/2�mS�L���դ�*��e#�5e�F�������t&��.�)`�e��c�"=5D�N!3,��p�R����
iK�(��Av[���u\H�1LHt+�{WC2�*RM��VJ�@�f�rE8P��	�