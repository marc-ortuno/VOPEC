BZh91AY&SY!��� 0_�Px��g߰����   P�we�s��P%S�'��OS&��444h@JA5O(z�� 1   ��B$�h=M4Ѡ4� �@i��&�&	��0`��$JdFF��	4��  dɐ� � S*�	>�~$Pw�&�_�d5�:��;$%P�)b�j�[��j���jlQ�؆��es�*N����VeE���Q�Gk(łэd�q����B�#ľ� ĸߣ���I��c�O�w�T����.�[������q��`I���,�v䖪FR� �*��jP�IUQȓiB�u[������K�^ @V $2t�-�[��Ğj$�KtފD��)*5i=
HP��aI�-S��S�聁���Η�[�����8b�L� �Z8�j�Wt����a]�ҝ3i�����(���SR8W�p�0!ZU�S.c�BJ�6(u����r���Y�Q$�n�fһ�q!of��VC.b�)�Z���d�t����F2�-c0�#�z����[<`E��'%M��s+�b9����<�ƅ2\Ʈ�d���u��d�@RH��IUr`�'�ƥ�⃩(�i}.E��)\��<�r�-� ���[��̭�R�^�4�E	��%�ur��b�n�r�$;����M���)^J�6�Ni(	�� 
%���@x�Է�(�(+�j��1B�F���>,3�1@�c\O���$A���F	�6��sX.@�PѺd2jU�č��g�/J���g�^ʔ#l�+BmG��۟A 5,��fˑ�U�L�L<�x$pل�(�Ʉ�zȈ����!,	�UPO�y.���ym$��O�Aj~�yUF8E�g���kk�̧W����ؘ4������"�(H�tm 