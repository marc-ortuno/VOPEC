BZh91AY&SY^֬� �_�Px��o߰����P���g 4!$�`
<"Bh�Q�&CM4 jzF �d ɑ�   ���T�A��b=@z���4����h`20110�L�L�	6�=4�M4� �47�!>��A$	($��Ht�,�[��F�p6� �ib��`a��Iÿ�8�����-z��S��#���N÷*Йa+��m��p�$]/�`Ή AKdW��K�L�$1�>N�ެ��T�`����#v1R�r��U(�\��fuHԣ�o�SB�G���-I��'pD��J����*� �R�5�ԡGIH ��D����Ր%�Yj��%43y�O�ԫ딳��Y��h��aN�scx6�� ��:���=��V*ǅ��N�)�0�T��0��XHb�˧Q� Fj��̥m�t��s����7#��GU��Wkލ��`���H}��oM:��V�"ΣW�M�}�h��|~"���Q�-��$l�'e��'�R��HP�Y�5n]�6�x���eר�&$Q�!�b�d��W��az69<�l�H���3ƓV��{��q+�?��8��"q��E�.�}����r�40?�C�M����a`e���
�xîw�1"4���.N*u,��95X�_���F{�JG���f��Қ�f$p�Sc�]�UGe�ڒ$��f�bG��x��sl9�MNP���Q�I �s�Or�R��I������01X�X�q�$YՇQ@)�o��!��P��$-�/e���a�j�8U��B�0��'dyVc&ޭ�HuH�Lk_N�#J$Y3�}#�jڅ-�	(�o>�ǖ{p`,���L,%@�+k1"������/�@�(5Ѡ)�|�PL?�A~X���/A��)��a�z�~����(OA�#%[ �X?�ܑN$��)�