BZh91AY&SYmi�< ߀Px��߰����P~t�&��I(��j��O2�& �Q�@h�F�hh�&MLL`��J��S�OH4�M @   �12dф�14�&��	2d�I��<��Q� OPi�b|�JbO��A�`M�����p�X�*b�j5[��r��i��[e84����Jpal&>��g`>��"$ǺE��2��	�ӤX̌��Q�@����?yCPƘ�um߭U�a9�M�I=P�p*����\eET��1ڣP����Nq/#K�y2U��XѕiW�C
BUI$
1�n�1�YF��&��y���t�&|��E1ND�.�d;����עטi�i�I%-��LtMaD��y!�Jg�ڱ�C����Ǣ��u,yc���SH�9�[F3ܼL�WE�K��2��v�ؠ:3��H1�Q!B�3��Ƹ�B�Q��1XL�A��<ꂃCQ���ܙ�nd��a�)�v��B:�	�����X�!��4�8�!�ev#�a�����^hT'�i���W�/���@P�F�|'m�#)i*�����Q%0�2`�����%jR�Stb�B��ռ�y��}k�Oi���L'�d(X�11k6�9�-�����Q�)$]9��|�^R�P&���$�8��&��*��3����P!L#OW ��ǌ��ܺq�a�o���jϑ@��bӋ��;5��UsNči�g��eD��r预j����eh��! ��_W�-�џ~���[zVLyG�bH�4>+KBѐ,
-��4%�C	 ���	
Pw_R��"ȴF�e��:|�7�,����rE8P�mi�<