BZh91AY&SY�b� _�Px��w߰����P^tF`QD$��AOA�$`F�h�LF���`&F F&&	�bi���BM4�����  hd�`&F F&&	�bi�� ��I��?SQ��)� 2��)|��	(P�D	?ԃ�`M���C^G�n�`�4��v�
�gټ�qk>N	���^Ѵ^��^N����v�FW�|��*'���Z��ș���`b�IS�����)��(r�ʽ��U�q�0ǤƘ�wժ��W��)2�<1���s둨�$\���2�ZtY~y��h�m[ɸV�!�!�:����vZ���D�In�H�SPE��R	С�B(��r�*t�i��a����a����1$w7�i�X5緙�S�Nfdҡ�ru^�k>ZHL0Zl;uXOb���
�Dw���&�hDw��NI��W�>�y�A}�����>&�����]�{��
!��K3��A���U��8���鴈�)Jڻ�VF�Nz9C *K��A;>��g!M5|Q�w2�#���,��bnT'��~�u�n3&%���xb�22!v\y�޳�$sҩ�A����^f�}D�#0����C�ӳ}n��(�U��)K!Ruqba`1�d�W�YS��D��s��2�J!@�S�2 �d�c�?�&�d�S�Ϝe�j�j�y@�0�]�D=�m=d��Z�C�]���ulP,S8������!; c���}Ie4�S��Qu)��=sP�SV�(�dA�a ������Uf{w�@V�~�k�*�Z�-�qn��e�ڵ7f5(��A�x��H0A� ��e�"Z`��	��҄���cd��2	mG�.�p�!r�5