BZh91AY&SYo�X j_�Px��g߰����   P�wd�9����J�٤G�S� h44 J�4
zjC��M      =D"���� 44�@i��&�&	��0`��$HI��!��I�2h4������1'�$!��%!'㓼��i-�m<&�<f�4����MV�Z���L���Q�Ԇ��Wȩ:-0E���|�?a31������I�A6T���V�c�aBRBJt.�$d\/�¬��
�1�>2�-��WB,4L-녀�3S�P�/�������j��$�(p�d��X�*�ܥ�I�3�4T�'������t��{0Ē��#�-��a�J.&�@�� HfN�{��l.��y���-�z)Jj��-R�Q�'a
��M�Ra9�E'cc�h�	 k�{��K㮘�ug˗���s(L�F���s};DF#�ف��;)z����9�i�_��*`i]Rw�GG�jO���/A�����Cb��X͏���H1�(�\�����>��g`�tf��+
!����Z���oT�y\>*��fN��:V�j�cKkH��5���RetZ���!M5�(�{�]��k1�10?�Z`�O���PxW�-��� (H��G�y-L�������Mc���X4'�ټ�D�I�0�f]_�k�4�{cԽw+UTߒaa���z9a1q08��+a���Q��H�9�N�k���
y^@L�t���j�N(8�W#CX����L#WN���r���G0?9��+�4WLҢa���n,@�=��(�$2D��*���?l��d�I(Q��A���J����T��i��U��t.���qO ����P���א�)7ǽmEúH2_j��"wK�#,"��!j�f1k*PE�!{��b		��*���)�~�r�