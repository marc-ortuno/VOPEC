BZh91AY&SY�B� �_�Px��o߰����   P�r)L�j�!$�&�'�c)�Mh� Ѡ2h�2b`b0#L1&L0i�e2��i�6��   CM 9�&& &#4���d�#���O��D���H��������F�`'� �������D�&K�!��#�n�bJ�H�KP��I�W�
��Aj��%L"�d���-B���!)
�B�|�2��`�v����j("�׸��:E���$��6HHX�g��>҅Ai���q��U���e��g��2aS�-�]���t��M��p��Ņu��d4��1P��{Cq�B�)h

���f,��V��.%��`Ad�+�XNw�Z`�z���jxbk��c��4lcco[m�hDe�o*x�i��;m�N�J)L�jT��2�I���p�r�0�]��� mj|�1~}��u}e�����S?����d�������3��L�i��gR�K��.��:�z�PD⪤�+�V��F�z;�Ns��B+�s0�U��f6���J�3��E����F��qpLF0�6)�=�
F���S��\�D@��1z�Xn�R�7��	 K�`��,"���˯G.�e� C����ӟ�Z��pey�� (H���x�0Dl!}D��a��]�x�xS�D�P�THN�4%�.���y�#K�6?B�دkND��m$�h�e
�F0�����0�	_~`jyK�"�I(
y� 	&N:C��K��}�.�h��q($B�G��A~���B�*�<��g��tWM��Y#��
3�]dvXb.`V�B4���P"d<B���)Ȯ~F��6�l(P=F���EW��2E���e5T�d��`�+����b���(�k8^U(&�A�܄��1A���ڬj�_�.[)��m'PE������FK�=��H�
 s�Y 