BZh91AY&SY�i�� ߀Px��w߰����P~t����J2zM4d6�!���FFLOH4�`20110�L�L���Ji�=M���j1$��0&&9�L�����a0CLM0$$ɑ�2����4���SOSL��	(P�D	?ԃ�`M��FC^'�n�`�EL]�C��}6���p��&�Y����Y*3���'˥��;�O�
�$�B�epX< ��"e���S=�B*/� �>ߝ5|
�4��V�J���~�䛠�Υ��#X2���
R��c�k��@�>$�LR����a�3�;�'�1������Ig�+~]���ԊCuoD�*T�O��U!3D�Lb�e!��T5F���ƛW?�Q{h~;���ؾ}^&�����I��V9MS��Nƿc!�1��������c.D��a8�S8.p-L ]��ؠ;����a��{�H^�K��[W���]�j1�r+
!��K°���j�{���f�"�*���K������/��9���!��4֘�!�ev#�������5�	��`���C]�����Q��E�.����4��;1�p .���-��*Gy#�˳
��ca�����X:���&4,�w������a��9��Fe�$��;���=e(� ���C"�!U�;�M��Q�E��t�:�S�۸C�OI!p�v�$���ua�㞥�l��{v��`�3��s5pU�;9&5�v��H�f�P�3U�l�n�H!@��<��UL�-�pi6���L�vL�^��<�Bѐ,
�4h
l�uC9 �hy�?%0Z�e�/�v���*�?�m.L./�w$S�	
&���