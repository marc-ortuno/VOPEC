BZh91AY&SY��i6 �߀Px��o߰����P�t
�f���"�	���"�����S�zCdcDmM4���L� �LL&4���(��hh�G��  � ��L� �LL&4��"A2S *=!���� &h�S��!P �H�'��>l	����!��7�
�H�sP��V~N+�F��fK�Og�m՗h Y� kCch?�����ft&T��q{Aq��{	˸W3f� �;$ ��}1��:	1�?�q�tU�s��O<.t�(�Q"��<���e��!�����ѓ�=�%J����FEmJ;��7RxZ�Ƭi&8�i�Z���R��R�^"�W]U���'u�Rn~s�cy6�����U��n�-�T2�be���d$�BL^�d;�aQ��'���6���!c����U�x�{o�Q7}2����"EBS���F+6�n]=���ːf;�EL�0���InR�>�����S��x�lP�!��%!D2mP����yw�~�gB�%�&�� ^�6��1PDWf8��Z�C
��s|l܊l^-���M.cF�
��k�!�����1&`����hoT'�9��=��\�L '#�ޏ��q�J�Z��y'�R����<�(�k���dlR;��g�-�Se͢\����\-U��'Β�b���W�s�6	�Vc�ήv�eM��	#9ϰ���Х(
x� 	&N:C����h�V}C0�X��u(
a��D=��	}d��5݉&'\����(6@����8��ubr�}*��N��S�ݼK�+3�:(GI�\(�dA�Q ������Y�o���᪙ԕd�y�P��=�C Z�+�Sx�iR�a�$k��Ab�!<�']�Ao��יr����V�,
�aw$S�	��`