BZh91AY&SY\��e �ߔPx��o߰����   P����M��J{SOP4'���M�h�@4h@����j@F��L	��0ɦ� ���4hl�FA�  ��� 挘� ���F	� �Dj�2dԞ�dL��@ h0�D�&�� �Xka
BM�o�y�؈�D	,l9��~l d18ؔ1���o���
""1�Q�����_5o9�MdH�i+�-ZQ�t��wQ�����M�c��..Ă%��KI��@%���B�i)!�L62���\tW96�N����%�a0�r��\ew=�q�K�4�d�ESD���8,�$�癶0�	M9�ܴ�14��(��F��|�X�L�p�EI�(U^�k�Ț@��0F_̄OSR�t���?)�DQ]�T�$��{�9&!7*�X�>�Sk��0A��#W��D��"�xe��$%���;��]��^w�49I�[�B7�Рu�>}�W��5mE�$�H�f�G�>�ݚ-�s�o�<�0�X��mC$��^��E����K	�	�*���'�RjO$�o����X��H�F��K`�d��R�fC'�R�ﳿ��y�C��XU�o�Ov-K0\�>nj�H���&4M�X�K&Qm��!��5���i��B��D��>Ӯ���C�:�$�n���Y#v5&{B��,�LT��G�����1�������z�T���
I��L�2:9O �\Gg aơ�.+5����]9��|��D 5�q��os���\����En�<d �Lo>��9	����$�ʬ��/�N,V�X/U@��v@ƌ&3O
�i!���0�_>bF��W�oiѺ�BVb"s1��$N5���]*~�m�gD��TJc���$MY�ww��дa�Ȁʕ��6�� L�I�mW������n#R���L����k2�1Q_MFK�02
W�1��.�p� ����