BZh91AY&SY��+ h߀Px��g߰����P�wd�8(WX$�OT�=D�E4cPh�4�4�@*aFJQ�      =D"�Ph4�C� d h��L`�a4� d�@�D�d&LS�3(� ���ğ8�@�P�AO��A�`M��d5�훀�"��T���0*jǻA�e|k�&��Cl{F�\�"��+HRt/��dfb}dr�HZ���KD�L�����б�B
�H0�`�(kƘ��kѭU|"ӄ���A��S:��pem+^)��r�B(B�1@]	�N�+�ő���Z*��7-Q�A*M�,�E�5��K):R���3x�DD@X $3'N�oZ܎�2y���.�)Jj�8�;��8�ЄHM	���&�Q�q�6� L�fw����k�B��;�|J�Jyn��7�z	Sa��g�Wǂ�WF���d�*��Ǫ	$Z�>�U�9��H��NI�Į�7)�A��[Ԧ([Y�2�\�hB�#�~ً�e�R�wX�u/OC�鯮m" �R�*�m�F5M�\���o��iX�5�i�FDɖZ�[L�\gT'�j�,@�ٔ.��L (K��I�0b"��KN�t�Y9�Ka0B�	6YV]"�3��(�>4��NFǩwޭUS<�L��#����nsp_Ei�1��$�S����ˊQ�0��B �d�c�?tL W���g�e�+�j��@P���H��.a����I�����%wӅdH�W6��,�����%EĆ�#"c\��%!�LӪj�j�B��"|d�`�\`�~�	!��5	�J��Yq�k�"Y�DDf�a# Y
�k�)�xn�Ge�qq�����SUnZ�2�$�?�&�%���Sz�w$S�	�A�