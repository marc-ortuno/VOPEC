BZh91AY&SYG��| 	_�Px��g߰����P��G9�P`Ȫ?T�4�MI��&FPh�jcRz��#C 4�� ����L&�@  z�9��& L&L  &M4$�J~�`�LLI�M��� 4�U����pH�@A'��!�`Y��L�l>�p:�3F��5���8v�]�n;��t��Z���u���j�X���}�_�߄K"P>�/Lܤi�b���
��.�	P] IT]��Mb���Yiı���`��ow���*�tj(N ��Z�4X�RP�`�
�K�֮n$��Т�|��cBH6]��5J���#%��� �0iRs"e�زkL���1DZ1�Uf�f�Ze\� .�Z��S���|���eZ<[��lccom��4�u��.��}D�V*�y��*��S�[�YDb2
�	�	���q��(����=�$Ђ�fJ�^�Ԯ�9��f^��,t�
�3�>~�EDnX���m���(�K�Ur ��a�@�j0lq�i��P���jt�:F��_x�L�:��)�k�1�H���>��	!�XP��R�����;�t٤HK��|�����.���^M?�H8�4)�N�-R쐛����TD��!3�d�G���+��m%�A�D<���L!=í���%֯�@ۅ	�������T^�z��+�'�J�L.:ofZ�R5K(&
LY1���8�[���*M�aA��
�dcp2���i)!��^W�&Zw��,��[��3�fte#X<$�'Q���!�����X�* ��p�a�ɧBqm��
�xf7(^���7�5��!5)��Zzr�I(QV��Fȩ�f&'8�N5F-��j���	�QQ��YA	HN��R'�;��YXV0⼐j���%��-���7� �삔� m���L�:���/D;�S�Ry B�ow$S�	i��