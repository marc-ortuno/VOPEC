BZh91AY&SYVd c_�Px��g߰����P�t��Ѯ�$�OSM4cP   � (S�SE<�OQ��    	L�b�CD�4ѓO�b4���L`�a4� d�@�D�����4ڍ 4��M-����\B}�D�	��h�C]�\�d��"�.v��SU��f��*7��XC���?i�g�"c��?���,�N�&]2�/'W��_�2�s��#2�	*TW H�:z�l���1�>�qkUd�XtL/���HUCb4&J
��冗���PY(�����`�F%���+�����@�%'��д����R70�rt��ݔ1Я5f:�BWI$
 c?^,jpx�hMU�̪`J�ҽ�i*�؁#"Hw"���)��rY�BQ��[�w�����^����m�:�đ�Y�>2	L�9㛃<.�$=��e d�h��"/���s ��.�;�/��a<���pR��nga��ƅ�G�1�g+
!�J0�@�l'6�{���3)D��kDB�M��C *%��A1kc�M5lQ�t2�۸��[�!�SJ�?1��W��^!��aB^~��S"3��Z���a������͎��#�H�2��_yL,1�f�Z�̬USL���#��y�Űݤ���6��F��Y�"��05<�۔��
x�0&F!`�K��<R��y,ڊ�
�0���B�s��$-��{I0�8_X{�tdP-�A�q�����@Ϟ�y�Z�iĎTƴti�%!�Lծj�j����L��Yr��zB�n���V_l����N��<D8��� XVqq4�&Z�!�� �HMA��������Q��"a���6+�0�*VS�.�p� ��<