BZh91AY&SY�qyJ 3߀Px��߰����P^rN#�	��*~�zR{hI�b��M#ѠM�L4hLL�i�      Jz����1A�F@��sLL�4a0LM0	�C`F"S�bD��#OI�@ 122]t��$%��V$��õ���Iw$�!��N�H`�(��jk'��nh�?$�+3	&�,mxYq��Q��^7+��Hٙ�n�"��JWŭb���~�FY�(Uy(��-�^_��;�
�WR@��Ơ �=s�a�PؒLi���y6*f�fy��SFӄԌ%!s�v2�,t��f����e;����HS���!����{�	X�P���(@�j���.*�&�����aa%���`�EdD�d���R�CCWi��Vl��EViY�E���1!_u��Yp��4��+�U �O��rL��K�b�y*©��k;q�n�I�H��$$@�v%��6���.Ƙ�� �M��E��;Mh(�郊��y�ӻ���BE��bh��W_�KOu��Q�#/����.�|PT��s�̳i6��'��K�s0�K����'�
 Ο�',�y�lą�$��_�@��0b�c��1�����s��t�DA�,���/Sٝ�B�U�5I��X�P��NJH�!�̲E���d&X��I'T�y�^�^M��LK	�AB\����x&$��r��ˎ
�G�e2`��PAcf��$����
=HJ�Ē��3�m©i��	��C�	%��9DŬ��q�3$;M����&ŉPe����[p'1�0��b �2P1��$��T�g �*+�j�94
@�|��k�bI~�K� �����%������r�G>���3@έ�~�d�jF�Ʒ����(U�s5p�B5�[�&�h��`T�y��������p`4/[�"�0a�)JS3���qp\2��j���zG~&&w@�`&�8���+S�9�k��b̽�(O����Ș5O�.�p�!��