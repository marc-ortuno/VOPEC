BZh91AY&SYe�� �ߔPx���߰����   Pz�8\hU/	$T𞚦�5O�M�4!�=D=F�b=55�j��S ��A�A��@1 �
h��i�ڐ�i�h ��(�A�ɓ&F�L�LH�A2zF��d��Hz�h��>7	�� @�H�'ӣ�D��4�P���Q���@��H���`Y�&G:� ��8%v8�;�Y�ˢon��>W<���ԍ9{�-���m����Tf�F�9B��_.��(Ɖ!$W�m��U=�ńi�U�����քf<��Ъt̍4�Q�k��X�*� $IULZ�j{%�BL��P!��8A# u6hz4�&���\L�"@���'C�:������(��u�$�gϧ���Fu��w�7��lccoCm�ilөk�v����&���M�]\K�X[m7�N͍L�C	4me'3�@C���l�	�&e�s�o.�h�������}5�wj���{���'
}$G�y�OoZ4�oƻ#�OS$R�vP��J�$�R�yx�����U��㙄��P8��D��)�I˄c��ص�M�[�ⰠW"*�6X.m�Q�e��q/�M" ���*�7^��KI����u�&���c$�`�i�g��;L�w�,`?�z('�k�,��Y�)i�a�TL��t�`a�:�=og�G�[!�{�LkB��~�ary�<�b�Ag�6��9m��6���Z5UG"��,��q�as�;a��p^Vj!�� �s�N��B!	8�#��p$���4;u<����
��Y"�vU�$LgQ��D�����F1�4o�m8\8������<�M�}jɤjF��-\2`���;6sT���(X3��!i@=8h�i��RҞQc�Y�xE���䬶Vl��.t� 1���9�J�e��6�	�� ��Qj�����9k����\���!��o�A��^���.�p� ˳�8