BZh91AY&SYRY#| �_�Px��߰����P�@fi�f��I$�4�Bx�'����1��昙2h�`��` ���SBh���=M�F�zA� ��h9�&L�0�&&��!�0# � ��ޒz�h�� 4hz�BȈM�'A Pu0�&���`%36�C��~%8s��3��t&�����p�I�q�v%��i��Cq}���n�(\��3�!PG�i�SC��;Q	zV��9ivD�tA{A	L� J������#1!�L7d�����tP��.��l2!��tʩ۳Ui�>�nT�T�Yؽ��+��z��zIk������r�y��kE��C�8���k�R�:!�K]j�L-f�!}Q���6r̙m��ʛ%���h������@��q�~.�x���(�"H����Q
lB��7����T��@����LoD�u��ptMͭt�2L�M��;�]���x�ܳ��
#^�{ٟ�d�9]�O!~��G�>c�A�����-�������Bt��O�'I��0��8��'�a���0���'[����_���[Ď�aՉXDJHs&p8�$2>��T��}ҙ�q�j�q��x�T:v,G6?��c 6�4S�L;.�+�Dt�,$V�D�{�jD|f}"���B���������L$;xr�D���~�4�3�L�z
����*���ƍA_q,hd$rSa��]�Nrؒ�`�� ��#�L.S����Dj�AQ��
��1�F�n�����_���{^@�n�G ��N��Xv��5�	�8H�M����Հ��i��+��J3�L���[�X��D�����z vH�lӣ�*���	�K���R�ѣR�ۦa�
�i���	�ea��a��+KBч�:UPKX�n�!0{�"���M�8�mC�Q���(���J̷�ǪC%R`Lg���)����