BZh91AY&SYGS�8 c߀Px��o߰����P�wd�;�uZ�[	�S�L��٩���i @�#Jy'��� �    %2D�@ddhi�   A��`&F F&&	�bi��!&
zf�z�O)�4 hOS��zĂ"��A	>=D�	��!���pf�i1nj5[��/�`qwY5d:��޳*Ӈ`ŉ<3��1���
���<.D�
�jM�
)��2&���0AD�F�C���ș��4��U[qUsB,<���yg�sH�R�:+��4\�*-=)ȩak
A��"Ӎ��EM�b��MJXBMh��a2*X�nY["��*���"������I�ϛ�cu��|u&���[SdʥISaf4�:�6(BHeBF4Rյ6@ ��h��i���E��CE3�чc��
CV�^�wQaP�ܧA%ߌ5��۽��Fy+�5J�e����OQbF�e8�W9��Q��� ؠk`�y����
$([Y�ϭr΅�G�����b(�.Q#������8r�7�� �3��+�Z�5�haRyr�HR�� f��n�k�+����̌��	��Ex=U�,+%Ĝ\���)��1"���6u]Ć퓦v���F��:��H�e�B���4�e��"��Uy�đ"b������q	��6���VB�IF,��|��ہJ!$�p`L"�B�]��g�|M��"Ԗ6���@P���b���x���I0�/�=�.��+��%��0V�3�y���S*C�"�ƴ��#*$U3f4P���v+D��(���������6	X_k�D"Bt����8����d1@�fL�MC�¢�a�$f�I(?Y	�T0EV��t[_%�j5Tei^�P)\��H�
�t� 