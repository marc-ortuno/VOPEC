BZh91AY&SY��� ߀Px��w߰����P~uI�$�I$�H{MI�h4ѐ4�hh�&d`bba0�!�&�	M
i���h�� ��0	����L&i��D�h�2LS��&�2�#@�5=C�_1>�%
-O�� �Xi/�׉�7�0UE�]�Cƪ��o�7����K?��6Uʙ�[IϵoЬ�˟%�(=�^��p�z�5�4S�W�Y��B��2��F��Tk�L���q`jX�]&B��(w���H�5}���Ֆ�|�r� ��6ce}	��0�BC�e�U];&��1��{m�L�6�ncW�$I��b�
j!B(S#�%!"+�2"Y���MD�ي�32���[�+�O/Y<۶y�Ȥ5f�����*1�hQ��R��Fƞ4�Zk��Ȟ�c=���-*o�Xq�]�pgz��=����!H/��Jb�ɟC^��34.����¡D3S�<*�6/o��>��M�DJY[3=8)�����/}|�6� C8�i�⌈#���ߤ��V�!�j7*���`uu�����	{:#���I�#2K}��ʪ�!~�
l �a�K%JC!�1Ma?��� \��a�V��@���r&

�
�!�&��cEq�0,6�bĒ0����\��	�<� 	&N:C��`y�T�g�ed[ՇR�
a{��{��=d���y&g\*F�*�D�ι��4���<f���ƶ��b��f�P�3U�(�TA٤�B��l{<�V3-�����=4��T	���(W�qf�@hȠo��B���U�Ü�h�R�qJ�GԦ-9W/��̵�O�EJ� �P��"�(Hi�r��