BZh91AY&SY�Қ� _�Px��w߰����P~tK&�h7	$�5=S6�4���= 4i� s �	������`���`%4B(b4�j� �   ��`&F F&&	�bi��!&	��bS���h��6D�l���(P�D	?������Ix���O���`�EL]�C��}{��7�����?����%,�*[*[���Xl>�sfH��E��`��^gȡ~¼��IS��@���}i���cLz������a�H	�1H�aсr���/;[78
�r��d��n���Mޅ���)���X����i$�3�|c��ݍK��"F�ۊD)L����UHC��Ԡ���ɦC�ʨj�z�z�W�u�������]~��q�R�0jkte2�a1rR�xgY����ַ5긭S8��w���ת��V��~;��g�����}�8�Aoz��Iu���j��څ�w#O�"����ZO
�F#=K���xf�I�ws�t���K&�	��^X	�GGM5lQ����q�ZL����05���"����
��G�w`�24��-�z��X�$q�R�@_D?�-eƕ#���e������"c�&a�.�*M4�H� E��t�Bae7���h�����1h$��= ��,
Q
�ytq
n��@`lE�*���9�S�۴CՎ����޻m$��9�Xz��gP.A��˦���-?�#>�\ӱ#�cZ���"����B:���(�Z ۜ�B��d���U3�^�Ui�=/��d��e
��\� X��f��<�TQ?y ��d �!.$�����m���:��`n�YX/�aw$S�	})��