BZh91AY&SY�-�� �߀Px��g߰����P�t�fi�H��@&A�I�	�� ��� 0��	��i� ɦ��i! Dz��2h�  4�0��	��i� ɦ�����FL�#	�@ h4�ji���X�@�� X$@����Xi.�&C]�l�t�V�"�]C�Z�5Z��|q��!�?=�j�(�Gx��!~͟�e�ݢ�*Kqu�\1��}�)��vs� ��������c�^�^5]�Eˮb��o�Y�[d�T/k\B��e7#Y�4fI�a%Fb��2�[fJ�Z��%����*&�e�RSVS��ut���E��O?$X�>�ȵi�Kn[A ��Qt��|�=�]U�Yw�b����5�L�B��!eN!XVM��
�P�V"Pw�I�M@�o�:v���e���K�5?r�B;m���%��\PlBw��_�k��v��P1����N�Hإ$�L�i\ޓ�>ȳc��ؠ:�#�2�R��H^bK��Ɲkp�h]B\��٤�(�o�KA�hPmpa�<D�9n�ڑK���sjv�k*
%u^k|d�ͣ� ���(�|̶�qq��,`��bp*�6u�0>t7
��Gd3�L$��r�.H��i�cD�����
G���fm�qMD�nɱ�^��ִ�$�0�@�%Ϡ�&�z�����0��#4�Oq�R�	�<r 	&N:C�D��b�Vr�Eb��P�6tk�`�KA �е\ `�8�-�U��Y;�I��a8`dm��]ƥ�$�$X�eWbW�&,tP��V�l�k�H!@�4�>�Y��Y��
�j�L�%@�+n��u�p�,��X�|jQ<d��C��`�ߴ�J"g���T���E'��fJ�A5��"�(HS��d 