BZh91AY&SY�܀� UߔPx��o߰����   P�we�;@���z2�=�= � h��d�h���J��S�ML���&� 4  ��SI��zF�@�  4 挘� ���F	� �$ �OFB`)1��#I�h6�#C$�>pA ��a�����]�"G{�%����훀�LAX�*b�j5c�ӿ�mD��P�<��Rg��Ĭ"o$�2���O�<���(Zb�"EJ��>�����g!*TY!�s�?mW�
 Ƙ�U���Y��S�\&�4�Iy��QX.�
�����UEʲAPY����Ee+B�A&�%L��ʊ�$�tU�Q�T]{�W{|�HBBJ�I L9�f&�v0�<ȑ6��R!Jd(��Hu�vB��"@!�"l�WTQ��17�(	D2��W�勎;��m��i�Q�,铫v$��j�<8q78'��L#�u�Y�
+��{B�2��k�D�T��7����րB��`.��(�)NJ$�.#>��p�H\��#?���B3���1Ѧ!�=tn���Lø�**�pʧ�(d	u��H&hk`Й�SMd�2s,�����^iT'�6u�(=6`�g&�
<�H�צ�B�Ik߶�+>�F�*L.�D�&:K��9#`̺��Zb�pl{W�2�uUMH$��1i u��(��t� �Ei�2�
1f$���`jw˅�(�@�S�9 I2p1�dL��\���d����("�6��!��<d��*�ra�ue�=;�s(����ǫP�A��gf�ͱY4ԍ�h�ȑT��͵(F�+r-D��`�g(�-K~�tѶ��EB.���
�3�̈́DF���ᐖ%k�)�|��Q�D�%�C�+��J�IL����X�;N--�L���1���"�(Hsn@C�