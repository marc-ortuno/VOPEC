BZh91AY&SY#v� h߀Px��o߰����P�t�DI"x���Ҟ��=F�M�4��CM`20110�L�L��M$h#@ �  `20110�L�L�B4��M'��Rz� ����M|D�"A+�$��B��V���k���"�Y���`Y��o�����~��ð���:��ښ6JL��Ϲ�����4�R�1+_�2Lg�ZL���IM��	C��t}�B������mp����ߛ麬e�aC�m0��`\�R̓�����E���E��G�u9%�AV��w�l����sk�j�j�v_8��A�W���� 2����_7�#}���h��lܚ̔�I5�,m��+]dBhB��Bc L�&�&E�a�_���wOއ��x��s2w����ݴz��2�$}�
Ѵ�u�U�Y��Fx��!�n��H�BM�+CS�Q�#�s0�ksb�D1'D'-�4�/��бԇ��H,alU�|l45����#��uiL��p;1U��������[�9:ETֈ�C�e�#˰�T���q��I^㗀�����¡%=���WNI��]�G_L�[7:��0��
Pf���i6�IC��w�����GF[J�kX֞	LX�#1W�{��v�=A�V`bX�K��Ƶ�W*vdL�&��@L�s񊁒�R������̐P����Cݳh�YAr�w�(���<��ʨN�8���:���;�.(�RU!��Ԙ��n��B�:9J�t�_�Ke胎��
�����͙��/�������$*R�*"K��!��F@�]pN���ġ�\H&~��q2�ޣ'r%�NZj��~��甹����K<��H�
b�� 