BZh91AY&SY%�� _�Px��߰����P^t�ɣZ1QO�OU=&�eFM����=@�� �9�&L�0�&&��!�0# �Њj�     49�&L�0�&&��!�0# � ��	�P�� �~�.���%
4�'��|i.�!������X4��w�
�c��ua�p��[uVz(l��YLj,Z�i�L?"�����BJ�l���-�^�&N]����T�������C�Ƙ�����WE�9��Pb��j��P�v��'�	%��9(���Ğ��U�iU���-z4>F��66�m�A�V�v1oB$�6�V!MQZ����B$F��l��єL�k�`!�5�^�m���B����N�:�0��3��Z�C�R-`����,4��G8�S�@B�{�:�F/��&aQ��>+��L��~���\d�d)ܔHP��g�t���F_�e�2�a�)�yUPbj4�z�8����q�J�\&;m:��:(G� '�!�4�4��FC��-G�iq3C�8�mT'�8{�=�f�2&%���w�L���.��4��H�Ω���5�F���jG���f�yL�@cj�!ӮX)�vɔ�XA`9� �kv�PcEi�6bĒ0����]��Q
��/2%�*:�y�]h�5�Z���s(���x��,Ϭ��`��$��s���8�Ҡ]w��y����M?^����Y4�H�Lkg��H�ήP�3VZl�o�H!@�5�ʬ�^��
�n�L*J�2V[2��Ȉ�w��� Y�th
m�U(�9 �-H��́ԗ�Ќ�DhH�
��{�Mh@l�rE8P�%��