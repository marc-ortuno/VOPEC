BZh91AY&SY.�� }_�Px��g߰����P�tR�i�BH�摒x)�1���#@6�4�&0a0�` 2i�a�AMI��� ��   s	�L �L&�  L�hH�@M4�M51&1�z�hi���)�i|�  
�J�D	?؃�`M���2�>sp3-EX��C�Z������a�(�/b���FӲ^�&�+d:?g��{8zaBeIj'[����f�E��,�I*T�!$`wΚ�@���n�䫔"�½�I����VP{(��g���E����Y�:$���v����T�$�2��~/�r�����Y�q;/���l5]�w�w�1w�_:2��������lx��]Ў<�!�<����bC��o��@J!� `0�&/&M2�U�����͈m6�Ht����G�I���ΞkՂ���v��/��ߨ��3�Y����vl�	F-�s��'U$$#bt+��*ˤ��p`��j��|����j$/Y%�g���3�0^�l�hZC6�Ka�j(0l�Sc�){݊0H)��h����|%�	�o�	��7@(9
i�⌇��nG����c��#r�?a��X��n���2aB^��|'�I�t�A�z�Qu�+[Lk��$7[��*G�H�3�o�M��6�ҽ5��Z�|��H����	��׸�tWA�SiF-d����R�ȥD	�>���'!��`d�R�:�Y"�T�(%
a}�=���<XfY��`�9f�4b�p���R�k�2{�F�*١;�9&5��p-h�Y�h�3V�l�p�H!@�4zzoUfzo�-����TƤ�%m�B�8�0�,�E�X�=YT�}d��!�$ ��Jf�1�]�n[+��}���x�d��2�C�]��B@��,