BZh91AY&SY�"ވ l_�Px��g߰����   P�t;�BI	�i=��h��4�2 �h T�eOSmS� 1  �  i�!MF�� M �4�ɓF�� �0F`$�!�=CQ��y4��4 =0S��I��ZlJBO��̉�
4���C^G|����V.���V���+kfV���96R�(�U<T�'��&���#�q�f��#Q8��\1�M;	�S�W���HIR��	�﻾�}e
�cL|j��9�q�\j��#�g#����uߺ�]l�������0j��Sh��	Ԣ�e_iP��)v� �JЦ0.��H� �ah���M&�,HZnI�� @V $3'N�����_�<�ID���%5R�(��R�RpM	��E&��Q�q�6+�����w�~t>*�Ȫ��M�Fx�y��Wzj��!��rj�6�{{�
�
��M�(�qe��.9bE��U�f�}���0�S���W���!H/�.�)��g��r���G�6~�K�lR��(0j5U|}�#�Gd�DA�lWq��:69C *K���A0-��L��W�G�-r<���,���Y��>��p����]�D�BG�ڏ�xkL��r�D��ٓ�W##�&
c@�����2#�Bޅ2��#}�6>��\:֙�0��Ѝ�;�N�1ss=���@i*rbĒ4�x�S�.�e(�@�S�" �d�c�?�LPX�T���e�-փ��(S��p�m��HV�\0~a�4d�I�ڥ��K.�p+duq=�
�Hw$t&5�ۘ�RRY��j(G=ׅ.D�oĠI@�����UY�>]h�o9q����L����+p""3��0	m(nѠ)�z�Ԣt�kC��0A��)��i�]�ZaK2����s+%k ��/��?�ܑN$5�� 