BZh91AY&SY�W�� v_�Px��o߰����P�wl�rh�N�H�鉒f�Tz� �h�OH#@h����=(f��@     )�M	���G�5=#6��4��`20110�L�L� �
m4ez� h���4���@���O�ȃ���Iq�k��7�bE�H����0*jǷQɓ�#`�3УG
j�uS�'�]d;F*%�Ul�p����}d�.y����JT�A����^��J�HI���dL�	�1�UV특��(�Rax�#xAa�S��j��̨�tt��^ak�Paz�$���k\�I+u����EZ��$f�F��+��_��
:�I7���&G�!		,I�͸�n>��M	�ĽSY�K	SZW�m��1��D�$�3�&�;\���kՍ��Y�C~�d&�f�$2��3��ڵ'\��@x<�\���Y���-z��}/R1M�"����`�8�<�|}�F�Cb��F��H1XԦ(\��fԸ�ԅ�z3}���)�p���=��{mʊ lvY[�������-8*O5�	�X�k�sP�Et�ɖ����P�����J�?)��YA�0]iya@�TO��i�r`�E�-��'7-=��l�&��� �p�ARy�<����Y%S�d�3�~_S�UTԉ&��H���t	�a�I�/�1�s�B�AF+�I��jwK��I&���$�8��&�/W����$W�F�N[ �<�h� \Cņ��t{񒙂�U�N�83���h`�3���e֬��#bcZ:t���y]|�(Fɫq-�P<F���ι1�j��.�kڷ`���6@�x����1��`P5�]aM#�uE�v2hD�� ��I�JR�O
ܾ+��k*RK�s}�Ę�:��]��BB�_��