BZh91AY&SY!	�� b߀Px��g߰����P����
:�$�M=#P~��= z����M �Q���LC�y@h    �$("����Q�&�S@�(� x��a0	�	��  	�M	$
m 
fAM4��4  @�Q'�H �X�A�߉�ZKx�F����j�ib�k�Iɟ!�h�q�Oۢ���������p���tu�z��v5ā!�t�q1�*�/��ص�IFE��C���/ j!�L7t��U+������g$��<�l���\�f�,�ldhT��j� E)e66,$��Q�Q+�%K-��@X�Bk:J�8> h�\�3W� �A/3m�i��<��˰�)R�:���lQ����-0��R*�b�ʦG��x(�hn( ���U��йc!.�����Ǧ�&���!�5�AA��KN�"��O����U~�
V)��3X�F��V��~:�?m�^9�Nu��k@R;�"���9W��T+V���&!��*h7b�ȝ��VNM�l�H����^u^}��,Sُe��8�D9�T�ifF��G%$��C:�5F���:0f^@�揜*�00�\9r�p�>�~C�Ih8+�[��eF	�y��y�8L�F���6��r�Ҕz�&b�F";zN�0���;�tT�!Y#",+���B�e_��1B&�q
&Vv��*
�T�5��j�DA9@�^����-+]t�`��6�X�-�8��ǟ@܂�@ǯyĳEDi����E�y(��r5��ab�8�`�rpԗ��`�#>�*TLak� ���'�)UƠ�*p�"��`G1��DP��z
���q:��O5��Q���'fZ��Wۈ���`d�g���)�O7�