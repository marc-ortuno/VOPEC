BZh91AY&SYn� ~ߔPx���߰����   P�wd��6E:�$�i�ة?I覍S��H�FG��ڞ�@J��A���h��  @$�#��4� h�4�hA��2b`b0#L1&L0H����4��M�Q�'��� i���f � D *	*�3 ����D��K�!�ên�bEcH����0*k"�H۱��������|�R��u�y1Jʟ3��%�\�92�Ml�K���L�=�T/d��Jt0��.Z�GUW�
cL|uw�n�V�D��Уx�1H�`h��[��\�
���TD���!R+-aFD�:��QiUƇy��Raл
L�����Ah4�Z���3�܎曬���Z�D�q������m�B�ޝ�β1dƘ�1��C2M�F�@�,�j��b�2iñʸaF�w<M��kqs�o�uC��9k�(nX��;6f{}�+�~���d1�Fk���ߨd��Ǘ�{��o<���
�X�z�2�Z��o
p`^����*�;m.�O
��=/@���K:�1z�Z�� !����fA��A��M魎(��r�R0X1�ڃL�d��6Q���Y�rA�'\��I��;�8��P�!��YA�x/��MzvVeL	ه.��>�(�+�<�k�p[B	7L����G���!Ȣ5�����ufU���I����4��b�8�6�VA���(Ł �9�N�q^R�"��I������0/W�r�љ$W�g1A(Sa�8�持t��u�`�6[ ݢy���.4n�=���gNÌͭd��#bc[�؂�*���R�p�YhQ��A���
�)�ǻR�Ͽ�2Eji�5�@��&yW�*�ߠP.	h(,����澢�a�$g�O���z
.T��Jn^��r"���Q��h`d��#/���)�w���