BZh91AY&SY�3A� jߔPx���߰����   P�wwwl�
�:�I�M=#S6�C@� ���F��ġ��4  ��  =E6��ښ �4 4h ���A�ɓ&F�L�LD�h�Sd�CCF��I��0LI�	E*������"Gs�%�!��i�7�0EcH����`TՏ�E^��2�v���z��\��ȭ:(�S�~����Lˏ��bG�Al��	%(R��?lt�P��$��C�"+Q�=!�����0���v�T(r-7L.�C��ͦNV�X.V� ��P��mF@�c����[T,�JwU5�xWA�8�>2�3^z�_4���Xۿ�k�(��K�����lDo�ȹ�7BS%3hۉ�*��&SN2R�B�q�2cL'-�.��A��.��05�ý����8rཷU�5p��ѽC���Y�D�"p�Va����e����8��|�V�y]w�n�ı#:�j2����w"[XG���`9�.QH0mQ$�r�f�~�jB�#�~��b(�gb�S}J�Q����8���M�DJUaV���g(d	tY��M��3`���d>VYj7�	��;�8�ҨO�k� zl�Ze&�
9w#�xnL�P9d���&�Ҭy��&���M������c1h;�f��"�s6=�ّZ:����&+J��Gɴ&�Kp�E1��+$aP=�<����(�@�S���$�8��&��.z��EqVm(
�6s�!�͜F��b�n^��f��r[]��c��H�f�\4�:xN3�d��)�h��#"$U3�^ʔ#�En �e����
����T��o�@Ff�[V#� >V@pΖUW:��
�`0[]aMC�uE��H0���
w��UY�5U�z�e��I/��FJ�A1<��5��"�(Hj�� 