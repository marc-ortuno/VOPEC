BZh91AY&SY���� ߀Px�ǿ�߰����P~t�&�p�IO�L�f�Q�CM@=&�C@� �0�M0  �4�0����44�  � � �0�M0  �4�0�!&&�h&���H@�d4�bz��(�"�wă���Iw����ٸ邬i1s�
����k���m���kޑ
��AŅ9���F���i�(Fi'��,�2��l�as9�*T_ Ahz;io���cL~S�j��D�3���M=��d9H�#�Ȋ&,*�]�T&�^pξL��J.@g�Ŝ{=e2jV����HIQ$�&q�{�� �"DH·b�
S!E(P���C1P�p�1���L�c�P��cw����Ν�t;�X��v�,:�E�wu7�����,�,ô�ǖ`�R�v��������:�[�YL���J֯I�.sk�F-l�Cb��V�ω��[�D��$���ϩx�B�s�7�9XQ��,�Mj�Q��������0�<�KSX۸������29-�-]�نm�V���؏&��f&�qy�P����+��0_a�0��.~���#)y%��T�Dc�5�pP�n8_'*Q��V���b�Գ�m��8�dI�b�?�&#~��2�Xn����EӞPjw�u�(�aOI�����"`^�R���b�TCU
)�l���a��˗E��x�.�=|�2(�pf1���x`�3�i�ɱW4�Hژ֎�&TH�f��P�Y��
6V�92P;L�?�R��g�pWU�����T	��ɔ+�""3�a�d���X��G���!���c��?a�4�J��Ț�k�ve��>Kf22X�����)��>0