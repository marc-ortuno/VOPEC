BZh91AY&SY�H?* iߔPx��g߰����   P�wd�:��HI"h��&F���4�4i�FM��0�Tħ�Jx�A�@�h  f��Dd�� @ �4�ɓF�� �0F`$�S��DѤ��4 4�M4hf���$!�JBO���;Xi.�������,EX�Z�Z��i-;�SX!��Uǩ.����$�P���*��+{�K���:�$5�V�R�MM]"F�!k!%J�$	���\6*!�1�tv��\y�o�4��5@P�c�Wl�y�+AA�U5����z�w؈�Ikre�Qԓ�T����	�y$ƩPx��Ğ�̭m-V�8�tD @\ P�{��<0�Sb�ٹ5�,��kV���I��sj��<b����x����wO����<b�^%n����{�J������ߎ����i�.��#�Z�k'߇��UT8���=Q[6LH��+��j��x�z$��?$6(U��{�q�6�KQ%�ga���3J��Y��P�����&N�5���w7ͤDJVһL�{��C (K�ޙ�S6�I�b�k4Q��L��w���0?�`kT'�8��]�C�I���&�t��"4[�s���p�;#Y
`���[yAby�<�f}AoiM7�ǵz�+�ZӂI��M�G���&�e� W1���aV=�`�xKv(�@�S� �d�c�>��,����2�D5a�(
�6�p�z��#�H[i\ӏ`�7S(|u�Rp��Ņ������ͅY)bHi�3L2��x���8�<�F��pSNf&C�8�Y zpԗ��8�ض�x�+�9�k�5%@�+n��+x���w��x�K"���X�{
�C�_�~��tq��Xg�]��_��f_��	7�ld��2	�d�,��.�p�!ؐ~T