BZh91AY&SY�� �߀Px��o߰����P>p� ;�6�6�I"zC�z����ꞡ�����4�@ h    )�#ҘjoT�i�� 0�h���h9�L�����a0CLM0
�L�)�Ҟ�)��C�z@ ɧ��N��W��Y$��H�$,������ԓ� ��y=w�˄f�)>Z�u�,��Ѝ��1�B @�c48~�$��3�ύchxZե)�6�LI+�Cm�5I���sNjb��M���g�-����V(�:Jz1�Ep�s\�n��M�i�(I1��!��z�Gqp�2a��~�&G"sTA'.w��.}��3Bi �G=�#�sGBn{P��i��:nC��A�D1�����B�ƣ��_[&E�&��2��+��D�uș�3���]e4R+,6%@YQ!�ug7��]mg �*�A���	j� `�%+&��kT�P�D��Yg'���^mXЋ��[3�ɇ�㒥�����4n:�1PBe��Q5������ma����8&K����+u��\�~to�N-o�w�ps�aL��X����Kıc�H �I�I(D �~x8�����;D��^Y�ʫ�עyR�l������m�UIt�T�#�BkB��h,�ݶ�P %�d��o��i9ɥɋ���������]��lL$���x ���jZ����"�6��3F���51�$Ֆ[5-X.�	wXH!��pq�E��SH��+��u?���\O��?n�e�h�DV����z�齘z)D�־7�;�����ej�le�i�ȼ�3����ԫ�Nkb���L��<{��3��$m\f��S��9�5ѽ�F�����u�RAm�+Ǭ�tGة�y��=��Vګ��Ry�=�N~�?�:R�8U+�{w��f:�e(��PGJA���t��|_	��Gy���b�{#���T��w�� �%�y�DS��+�;@܍Ȭ�F2`ڋ����r���0���Ā�-/�!�g5e�cN�T@��pk@��Iy�:�$�:Eʕ:�~)��?�9v얎��9�U4K;5H8b�5-]������X_h�M��6
8� �>ŭkt�n7)d�0r�n�UѮ��~H��lA��:T�D����d��R�]���W&A=��ܑN$��@