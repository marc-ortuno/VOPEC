BZh91AY&SY�Ë ߀Px��o߰����`<x�� .�@4�	$�O@���M��z�@b��i�S��4�� ���  44 ��4�   S*O"�yCOSj 4 � �`&F F&&	�bi�T�ii0MM2i�2 h���bj�@�"I!	�҈,���՟�ԓ�KT�x^�{�H2T���5-�&�x� �!@�1��1�`�!�lc!�M1��1B61�B1��I�a�:��ٸ��p pa���! Z���dRi2�)A8����&arAI��m��MSe�	(�C�h�w�����v��yY���6+��xzSSe7�#��g��X.�@R�+�ߧ>ɣe���]���6�L"d�bR��;��xC}��#U=�к;0���$WW�,�o#2@k�u�YG
,�U�8+W�+�̦����-m-�<@�_�c���ԭm!4�J(�Vtv�Z%Jݢ�@��6f�Ӏ��WJ�d�
)�uw�V�t���ޢ�:��_��3�����%�h\�"��"CJ��b�&�	��*A����=���ǭ��T"�[�r�����m��w)�j�*��qP�U5���3I���QIR1eH�\����7@�FoWo��'$5��9"�M�|yR�Vn���8)g/.�ܹ�[�4)ê{�R-6J:�A ���@��!��GqgjH����ˮYiD���T�V
s+7��͚5s&��ˉt��|��0�c��G2|#�$H$��$�j�  ������ja
����v^#fX2�4*!���	P���А�%�.	R�SƗ�jΰ�b�cS��\���H�ͭΕ�s;�,9H�<�wWҡ/��{z�a� L [Y���f)�]zl���T����X����Q$ ^�}W+����� 5-T�=3S�������w�.����8tO:"z����d]$cm�����1R��8�ƛܧ~��:���� "X�*pL�ٟ��eP�ԩ�ү-5[Z��2�8���LYP��*�\�+��^��W,�snd��п��~�ӶQHnZw0�=�x��;o�~)#q�?Mn���Nns/{��:s�T����3V��I#	Fn5(g��%'c���7b��yNf�;M�k�qR�p��c�H,�c�ް�R�R��~6����7K駙L�i��hw� Z\v>\B�j�@,s.I?��D��a8[����ǿ�]���=���Ω��g#�R�?���H`�quu薎����3K:v����n���XT�wˬ�s(�^EY� ��Zַmf�,�؝Y��c�[6�b�7�0 j'gJ���ɜ����Y��J���dd�L�9��.�p�!��