BZh91AY&SY$� h߀Px��o߰����P�Թ��tDI
~�x��)��S�h44� �i�i��� ���	���OP�Ѡ  ���L� �LL&4��"AS��LF�!�6�T�Sj  ��=M2�$�Ă"��D$�{�20&�X�2�>pSX4��x5
�c塾���XZ��(���ùF�i�D����}��7P�RZ�ŶAh�^�$]��5��HIR��F���S_���Cc��������0��
�����cl4ja/T��R�.Q�qֲ��h������!&4���g���Ol �.x�,賉aE Ѫ�i*�<l,���5��/$m��lDyi�s�p�E	L��k�e':r����2���fBc$Ɉb�ɦC�h�
Q�e��B����*���.Z��+���]�N���t7�2����2C;+�B��Z(�Nx�lB̈́֘�"5S��,Y�x!�XG��a88V�{�c��sQ!B�g��E�3D.b=Q��`LE��S�|X��,.#޼iR���ש�����/>R	�k\	�E4��FC�e���.&u0?�07*�8x��{��0�Ę@P���?)��0b#a�%���:,v�;r�a��f���j2R=�/�z��1�ɱ�^���i�D��m�G��=�b�9n=���Ӹ/*m(Ű�/��S�]��aO�$$���H�L
Ug�gT��5S�@P�ßX���|ą���q&�tJm���];���c�6�T���qKC�#�1���؉���#�Ֆ�,Dz�(�o?]Y�z^@V�Mt���%e�Bβ"#=F��2�@�oWPSp��R�a�$հ��N�5��'�9B�-6N̾�ԏ�1{%s �����"�(H��R 