BZh91AY&SY��q^ h߀Px��g߰����P�t�II�jz��oM$6�G���� hh�` &	�  &���E h�� �0��	��i� ɦ���К�OScJhhh�O(ژLI��W I�~��m%�!�י��"�H�sP��V}{�:Z��� ���^���RI�B6���RO�_č{�L�h�R2'���%���]����RBJ�+ H�=�*h�
B��{3�U���i�
m�36<XnW��rv��$]��̉J�	�Y�!��MEh]�)�1����q�0�F��2fm,/�Wh,�Q;��������`Cj/��5�Ģ�lSb�7f�%�RMkAc&�b���P�H����V1A�M����x����/�1���+������|�Pv|m�<ć�z�0��r�4Fu
�����{�����iU�˕�&�w��G�rN�T�nR��R��rg��z���G���}���f�)k<����{\G��	���)Jڻ�f�*r��R^��d��0L��XEGk-z?�a�2���Mʄ�����{��i��L (K�����Ҙ1���Iq��Oz״��:��o�=��#đ�f;ޅ5�f#�d�65�
��P�W�I�1�D´Ɉ�TW��ASiF-D��s�OL�i)D"��I�����(�@Z��;��2�.�j�2��L#�����=�;I�B���S����nJ�316s�>���3���2�V�C�#�1���jIHefq蚄t�Z�e��(ǳ�U��o��������%k�"��11F@��7�pSp��R�a�$�Y�qJ����S����Y��Z|<bdd��j����)��[��