BZh91AY&SY�� }߀Px��o߰����P�t��ɦ�!$��h��<jG�h4 z�P�h� ������� � A�@  i��ST�C# dj  @ �0# #	��14�H�S�M�OjC�Tz@=@��jyOSԺ`x�A%�O�� �Xi/0L����)�"�]�C�X�n:0��]��2�B���kB^��읆L�?g�7���2��'���z�O�V�3$��MRE���L?��Li�Ҷ�⫌"Ӝ¶�^GFR0��� @�pV��,,3p�L�!�-�u+H�: $�nܚ8@��X1�J��Bb��6�0���m�Q(@QIRN����66����[�.�GdP(
��R��T�|��������&/6M8v�VQ�����m`�ȋ���]D�����e��V���ХyYH)�H�-�+�%��c��u��8��B�zJ����Õe��wpB�Ć�֮9>�,� ��D��g�׽y�܅��:�`��f�<��QA�Q�[�!w���,��=)5�#֌W�r�(����'�Nj�FC�e��˨�����q��P��p�� {l��dL (K��	ߊ`�;Xr��Ɏn5T��+�0G�Jd6��H����0�z�i�.�u�>+�R�u�7!I1Zf�F`��Q�&.������:��Z���jx˫�I&�Ȁ$�8��&+*��3D��5S�A(S�ۼCٖ�_I!p�v\I�����J�t���>{��2h��ux+&��H�Lkgn�Z�"�:8QB8�YhQ��A�I �����U���
�n�L*J�2V[0T,�C����d"��n�M�ӍJ	���_��?Ă���-�s��Ԣ̾�����d�X:��rE8P���