BZh91AY&SYQ h߀Px��o߰����P�t�DI)�#�)�3SCM�A��4ѣM`20110�L�L��M(�4� h  2 �0# #	��14�H�F��И�$�z@ dbyM4�bO�H B(	\ �'��H?��K�C!�#�7�"�U���`U��_�_Q��a��a1�m
�h�Q�7�_Ğ���hL�,�ů���2�LƝ����䄕*k�$b?
a��9�cL}^wl櫮c�a�|(�|�3G��l�P�/ib��+}�����89a{�V���'u�d��&U��.�;��n��������YO��Y�[K�I���:�"!4�Ύ�p�xS�M�m��Y��)&��X�ف�PM�R)P��H2I��Ȱ�7K��bn�����W�d[�s{-]�׾f�Va�b!k����]z)��Q�(�V������.H="���ıt��_a#���ƥ8[!E�%ȝ ����}�b�,�6"�^FF0�F)�>5
F�����v]�6�E)[����O�k�2��o�H&��r&s�XEɗ��Q�2��!�f�B~���Y�~����aB]��3�4���d.�K�O:x-��;j�c�
�4~�7��T�G!�n�Jm���6������aִ��$�cF�h#��;��:����Ec�2*n(Ŭ�2���S�]Y��aO�� �d�c�?�&k5*��2��j��@P�˻�Cݳh����d�p$���<a�WS�d�LS�����@Ǎ�����=	�n��#Z$VgTP�sW�(�z ��H!@�4z|�*�f�2�+��U2�*�_i��A�&!����\�=YԢ6��j7P�É�g�CB��Ȓ���U32�=C�Y+���.�p� �$8