BZh91AY&SY"�c~ �߀Px���߰����P�q#��0�I%6��&�4Ě=� �@h �<h�M@�@     JdBL�z�P��� @�4�ɓF�� �0F`$�dhL ���OP�@S��b]0B{ �I��I��$f�K�d5��񘄬EX�Z��d�o��|">��!��1��!�biF�q5�vS��em�r�t4ˤ�E)m�ӅR&�%	˪����uv���v(�+�ŶAh�e/ę��B���I *Y!.�
]��9@c�=���B&vL/�U1fe��CU"[yxI���"Գ�cn�%q!���1�h�_5VxV>�j�!D`f�fɳ�v���r&`Λ�jI�"�b��dh,�E	$5v���̮	��BШ�* [�(��c ��V|�)D��M^R�L����BE 16i���AwEP�Hy�8Cu�ӵg��L�Mp%��� 0+'�Q@��������4�N����E	Q4wׂo2�ĩ��BxmD�8!��	qH(  �t"КԦ�(���23+��Ε�s;�=�b8]����h՞mm��Ҵ 8�q��G�U���B�Ӄdv�%��]�Oר��Z�
2,���y0��s0�U�C�h�)��1B����Z�3���F?���"��)�:��5�v����3iR����>pW�sb�R]���&7Z�Q�Nj�FC\Yd�Q��,`z '�	��ݢ��1-3�	I�����L �9���;��F�G65L2�Q��Ӭ�b�v�7ͨ,�)�����[��Z:֜�E��!C$%@��2	�YeF�^y��1��Q�9 �9�����)D��L)렀&LB�^�@B6FȬ#�FRa�8�)�o��!��H�	~e�q&�fk������W�J9p`N���XM��� �D���׬g@H�2Pݾ��5m�F�E�	(Ƨ��b��V��dn6_L�%@����
e�H��9L��dA@�nL�Mc�
��H�4�Dه��X���D�R��L��쾟R2U�A%���"�(Hz�� 