BZh91AY&SY߲D� _�Px��o߰����   P~pS�#rhЪA%
���eC`�O(��@h� d����
       )��i�=OL�M= �4�   �=@hɉ�	���0 �`�0�BL��OI�S�ɽI�M4��jz�C=D9�FE� ��� �>}����-
���y�X��T3�ȍ��0Z��?b�1�!��C��C!C�<Ǝ���)�_9�X[Z�+$�I���3U%J���!J�J�&��t����l��;��I���b������]�er����29& �8� ����v�qb�P�#����ݔ���ŵƉ�]0�ۗΜ�ISES����-E�ͦ�L�Y�*�;`�9oXU\�$��@2r[��'2��ba��{�2�Ќvأ%�ؚ�2��SN.�j qA6�ւWа�LJkN#MlP��R��\��(b%ܳh�'(�)�ƛ1F��-E��)b(6S�ѸRu�A̐F�}�4Fl^%���m�ٱ#Q/z�P�r϶�N�Ӗ`�HN��W�͚]�
�A1SN��`P��+1-�K�y�L�̶�[��}�A�ԙ�j�&�2$�h��v�6@��G4�A!%ĒHD@1��u�S��h�MGqwf�*�J�܃zFCP�2!� Ƞb��)A@ �ފ��*n����.U�D"����>�����_��}��-O����#�.�d 8I8�c[��O��Z���r�v�Jߜ�O��uB2^R�$�fU_׹]��nP��	 ��2w9��Z����y4���A�k�����k�v�El�c]G��,�����M���J lv��/�tq��ݞ���'Ǐ��U���tU�<�	���`��L����D�nlW�8~���a�E咁qS��ڹ�` T'"^�����޷V҇N�Ɂ�I�(e�T@�8�aF���|�	!��\A�'.���h�`l��*���`|�V�2�R08��1��EMk�C\i��AIx�$
0VH"�٨��95�|��P�fǤ�KP�/.F��E �p���sI�7ê�uSE���(�X�A����u�����,��T2P��H��j�Qk�����i��l�ɣ"V���WF��1K�.�p��n)`�%/�¡V��fgv�@h ��X6a�0[y��X`;4B5b1�Am��)��KVz`�-��y�bbV&JFO�z?�ܑN$7�8�