BZh91AY&SY3��[ T߀Px��g߰����P�we��L�u��)�d=4�����hTi��
##A�@ 4h  d�MQ�~��ڀ�4h  � s	�L �L&�  L�hH��M=54��h�=56� �b]0O8 �AA
�}�2�m%�C\ٸ��,EL^���SV=����l�a�b���C�� w��XGڻ��WԪ�¤���B��)U�B�ːs�9�/��\�i����4���eڕW�-7L)�L��LPm&���X.�z�L��
58J@�:�`=��fu����g�I@JE�i�UX�~���P��i�5�	:�@,{݅�&�!�w�n�P��>J�Q�R��W�pe!��Hj�z���̪mnu-�����O5��c�u���^����@q��;w�.�K��sơ�R��iz���~��h�-�+�y�DW��ڡ(�q��0�R��Jb����*�32�<���XC/b�}�@�,�6��)f��0H(��w@
�m�D TK}�R	��HЙ�SM]dA�e��s�,`x���*�>�O`��g _i�0��.>Twܦ�``�r���L�1�*`��
�%vH'���#�'�I

�ܢ�n��
����d�Zdi@7��Bb�s�6:+Ma���(Ō�1Nx���-w��AaO,I�����0<DcX��g@�$W�F�!L"�L"j���x��e�=���pϊ����K��L���0h��l8��&�ڑ̘�/^P1�HeS4i��j��Уe��? ����x�U<����$��u�
BSP������B� X�XS(�諸l�,/C��q �i$�NE����Y�µ$�t̖&AES��"�(H��-�