BZh91AY&SY!�2� iߔPx��o߰����   P�wwg昒�	$L���=Oh��?Rz���=@C���Tɔ��M4�      S()��F�� � �4d���`F�b0L�`�!	�~���S&M�� 4 d�C��I��V�X���f_�?L
4�h�C]�\�d��"�/P����>��wԂ���D�a�J/yK
�����P�O��~�d�>2���2�jPMu0b���(R�$�/�����6{H�&8�;�J6��»�&4�#qRÖ�[h��4���7�%���.ϔ2i%�I��qǆB�Hͪ�idU'I�^�[4��8����9����d�
n�����H@�{���=�Д�L�[R���BJU�To�&�iQ5 DcD�5mJ�
(�qf(H���n���x��	e��>9��*����kۍ�$�A�)=VZ������Vss6�8���q+��N���;�rݼ�;���;HlP�w��H/ڢIB��ϩ~FiB�#�0��.	��A��x�T��+������56:R��`���Ri�B\Vx�&g��1'�'5
��!��vDo�/&Z��!�LU	�N�Y��vp�Ch��#g�>��T���G,ǭym�J�y��L~�A��<
����̓�9�D�k���m\-R1������1{��X��t�R;�Y�+G�s�5:˚�(�@�S�� I2p1�LL
��m���H�!�M�B�G&�b9��<[k^M#�;���o�8YT��}Z��v@ǳ#2͋E	$�����"�<��fا#,��2
Z��(P<�/ՏF:ꋠ,���a#:1�<�S2�B�b1RV�4����e¢~��:yJ`�3B2h���}Lˑr�?9�X�2	��.��]��B@����