BZh91AY&SY�&� �߀Px��g߰����PXypmrd�	$�4��Q��� =@=A�h�j`��       	H��z#�Sj==@  bi�C�L`�a4� d�@�D��i����� �44P$=���@!,�	>�K�K�2�9i�sЁf4�1xچ���;zw ��-\Ns9\?��y�����8"`�qTʒb
�������M�`��qepX=�\e��m�"���䐑J��!����,�� !�1��b��U�a�0�\)���٭�D܍2��	7e�z'!��[- ��+I�+�Y��5�[�AI�������0!5�Y!(Ȩ EeI*&*
�3@�T0�Z����d{2��:X��!ł��#�����z(49GV�,��4���	��lTr�
�oÑV ��XC�h�\�;�Heɓ������Ͷ��DxjܺadP�ɣ��'.��8�l]���d
` a$�Y4���Q�NG{  fT7Ӝ���wT��Ɏ~.z�TF����˴H51�y���6�KF}��58��X,e�_	Hؽ>��Xo[��8�-�xؠ:�3����)>�)%���א�h]�#�����lS���0j7���G�-��"��x�mҫ���8E��ϪB�K[]р>!:P�E��+�[�d�L�qq�P�9��V��^p���aB]a�<�&Fb%�����~�Gz��� ��a��gR;IF[�+�)�� ����̬UST�@�ܧ8��N=' f����
1f$�y���-��@�L/��@�P1�?|P�}N�fRU�GQA�0����z/�9Im�~2L5��Jy�Ĝ+^� �[�
Y���)a@�bG
cZ:t��ȑT͛h�U�l�Pk�H!@�<<�*��j�+���--��d��`"�zȈ�2@�2y@�f,AM#�tdB`�ӌM�p��"�HP�MUn_���j2(��b�J�A5��"�(Hd�wM�