BZh91AY&SY�J�� kߔPx��o߰����   P�u���i�"H����m$f��OP�'� zF�i�@�lAL�2     z�D��z�hh��  44 挘� ���F	� �$ #M�'�M` ��F��=� ��%XM�HI���"G�F���k�ꛀ�"��T���0*j��^��2�v���<�k<�d�`�'D�l���{{�ӻ]�&TKI8��-�^_��Ir
�K0zP�s�"������@��0���w~���M=煭�i�g9��.6�~Y�9���9�[�����@���B��RQvP��]�N�I��P-�F ������D�68���p������`C2t��͖��𧚉(��7b����Q��S�TP�BhL��E&�����Llv�`H���l��|u����ygO�f8����ߣ3vi���f0��Q����Ym����/V���+h�QQ�G9gܷu�|�F,#"��|�8�Aw*�%!�����3j(��c��XF0�c�:�
F��G2��yΕ�X�.4��q:SQ��JL�Ot`��)���2s,������`d�O���@<��ZbM$q�#�;�L�\9m�e�=F̯�`��
&�9�+/O:��,�)�!|���+ن�p�Hh��L)d"b:wA0�t��t�`����Ѣs�O	p`R�D	�?���'!����`��\#,�\CU��B�F�6bZ��<Xؼ�`�7�Hpم��ʷ����78hd{�6��T�Hi$d�e��H���9��b���+n
6Z�73�Q@���2yw�f̳�@Uq��h��d��b(��""2��/	l(-�����¢�a�����Az����O.�+f]��}dmd�02	Q�/��]��BC}*�4