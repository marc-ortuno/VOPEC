BZh91AY&SYf��� �_�Px��g߰����   P�t]��
(BI$cS$�i����F��F��
�?AM 4h &�  4��j�@�� �i�� i��&�&	��0`��$H &Mɔ��3S�@ c
mB��@�@�� X1���y<�i/&C^'�n�0�H�cP��T;���Y��m���3�������88Mn�$	J%���y��&T�I���p��j5l(c�`�3e�@*V@�����(TI�1�U�y�U�q�e�
C�Ub��N����k|8��ʻ�]-I;=5"JN�-'
��M�*Mf� ��G!iP��6 ��@%KX0�\S�L��)�o���*���e3�861���m�i'=������R�M#(��AT�8�ɍBc����d�!��d5F��C2��Ι�4;4��%�r�%r�V^���D��g-+�n�Ӧ�}��O8⒢�D$���TJĎ!	��4�	-Jэc�>ݥ`a-��88բ�s�(��@;T��.��&��f�.�/�4���̘���(��UW���xY�6�E)[J�=Y�jT磔2������Z�#ΑM5|Q�y�ۑ��/&Z���8�ܨO�q��=��\k&�
=���g�I���]D�}4����zU0�h4N�K�jG���f�𦻍�>�a���'�va`y[ U�e�q	��a���\sJ�J1fI�y�S�\�)D
��I�����(�pk5>�`�t�b��(
a�x�{�m��,W�y&�I����Ӆ�g�6 ��1ل�-�R�I;�9�5��p�i�Vg�Ǧ�ʊ��"��P$�x���N
�ٻ�H���3�5%@�+n���H���!-�e�X�=YT�u��C��0A��)�Xc�f�^pmy�+2y<�d�02���U_���)�4}O�