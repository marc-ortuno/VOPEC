BZh91AY&SY�ℳ iߔPx���߰����   P�wd�8(��)�LSi���b� �4 ��T�SBhzA�  hd  ��G��i�� 4�   9�&& &#4���d�#�&�MO�
�����Jz�� 02�yCDĞ� ��%XjbR+�R$|�i/��O���`�ƑS��`TՏ���i�[F����Hk�Q��`�'D�����{}�ʹ���H[��&����b��B��_�T��@��o}�
�{
cL|��V�N����۲U���Tf}��Ѿ�V��jz�����(�­$pbr\�aT��.��3B$(��zl���+2ڱc��Q�G�/�|�D�!�:u�sp;+�I�J$�ؤA)�"�eD��`��N���I��E&�"���Ll6@�h�w���|5ӑWU���*�+�����ޚT3�-P�U��y�����l~��HJ��'�U9bF�d�򬹏�x�L#JrN���1�R�JiB�3�׽c7!f#�����e�R��Pbj5T����
�H�"��­�<jT��"�_u����p�����(Ȃ;Ye���h&X����j�>Ӈ�- �٬/�Ě (H��t�0b#BJ91I�`�y��SVە�N`O8Ǒ�M�SMb7ۋc�x+GUT�$��&�d#���&.ÞӠaEi�4�
1`H4�xS�\�)D"x��'!�Q0<�`�S�YQ�Ȳ!����0�>���$.:Wנ�3�M���R�s�e�]ۇ�1h��}&�
ɤ;R9&5�=�0IHeS?��P�4V�
3��Z3�HN�ȩ[#}8%��RS)*�Yl�QY�qm��p�K"�����=W�PL:���'�\���SY�n[!xl���+R]���c`d�n���rE8P��ℳ