BZh91AY&SY^&�@ ߀Px��߰����P^t�f�h�II����f�)���L�Lh22U��z����@ 4d  JhB!4�l�L�S4L �&MLL`��H���h�!F���I��M2&'�$�A@G �}���	��p�k����v�cH����`T�o	�,k!_���~���6U�I�8�Կ����S�&
T�$ŕ�`��̰&[��+K�)$�:� -��^�1�*�ϹU�a�0�	�1H�aB�cB��.	�־��L��"����Χ�X���7_�D���לF�BXIg�ʹ�.ƾ��D�&�ފ�)�
_XH�"	��%���Q��U76�L�ʛ�����d��$yi�l&���Wj|7��/��xkk|UBƍ���	�_^�
a���s�7<�i43���в��� Ɋ�
�~�8�p�,O_���)A��y�R(��f�u��?V��fǥ+us�4��(t�P�k��5hk�am���(�}��wr	�ф\jT'�l�(=U�X^L (K��?���������Ƕ����8�0����F��#���f]!_���0�Y�PqV*}�EP�Aa��]�7�9C=� e*4�b�H2�y���.K�Q
AOl���q
��/ clmF؋AWt�1(����C�~���e]	0��=;t�P-���i���{��m���bF�ƴ��3�ES5좄m����eb��1 ��hi��ǟM*h`*��8X�.E��DId2F@�(���
jk�(&� ����D�2P\�J��q���!��Z��&� ��?��H�
��� 