BZh91AY&SY91�� �߀Px��g߰����P�t��YM�XH��J~	=S�MCM�yG��C&�����` &	�  &��P	M�yOSG�zj    s	�L �L&�  L�hH�Q�M5=	�f��h �f& |�B��H�'�� �0&�\D�q:��;f�4��t5
����u��3pv�ΝS?�Cn�ƪ�j����O"c��q��<v�m�2��'e���A�zI��yEi{1� )S	 +���K��Ę�uspޫ|#����y�oUɅd"�)����f��n[�1��fq,�r�I4T��2�Tˏ7(kAV�!)*4���g��H�t�tFLqe��R{t����$�&fqϾ�[��Ð�"H����Q
lB�R(w��Y"G3$�&$�ŔL�c�`!�5���ЛU>0�W��L��'��N��(���p��R�L�G�����!)԰�m뫆���f�.����j�%ei.�\���>��ț%�A�@:'��,�Q
v(D\�W+<��_��!l֋x\N!��FӍ�a����qN����fǵ���k�Ogj�C��wO��{#H��&�������G.��fF�I��B|�"����}�����t|�m��-��m���4�9�*��Q/���R�i@ʯ	��[Ap�����Z�r֚�Xb�,D�|G1x��h�����J1h$��= ��=�(�@�S� �d�B��K�cE#QAN��X�A�w���/qh�k��C�T�Ӧ���,L��A�Ɓ��5�)�$�	�5Fq*�Y�6�B7Me�(ٕr�$�y�^?�j��y����KgDX$������yA��e�25=�(��An��Z�ݸ��b�"����+k�j�o���,
*��.�p� rcO