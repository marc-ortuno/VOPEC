BZh91AY&SY3��� �_�px��߰����P�p��J�9l����I�G���)�hш��24�� �� � 1   HDSOTm��=���M Ɉ�hɉ�	���0 �`�0��$)�hMI��F�yOP 螓C[��,$�)dH�I^��g�B��y���O7��c�zH�*F4�V�-h�|Μ<���0��d �B"bjd�@� � ���W�ǹL:\�Z�ݩ���t&���Iu�%�W��ڦ�+�?����C��q�fWh���fj�,�8�k�ޚ�iu�D/���Y�ya��`�!)R�������h���Ƭ�َ����Lxæ�WMGW���m������˥w.fƘ]�
��f~f���ɋ�ǳ�e�k�S��^v"�mԣ/i,���ᾑ�T̼Ecw��n�9�!4�1��;�a���r3V��ť,b:IL�93��rFj��Jc$1Ut^'��ٝ@����eJ�hp�ZwP���T�$��k:-�q�ZtD��T���|4Z�*�J���7:������̻�ie��qL^���r1L�&�A}�G@j����]�2���j��#�l����U�Up�Z��O�sf`�M��M����Ո��bF껁,a`�tѩ�k������l(C�����#���*ʳ��*�S��9��a7D# @Ɓ6ٹ��bHbC;Y����`Fe�Cf@�̫��:��٥�,�չ�eQ�X�����I������o O<���YtѬ��� ������Kԥ� Z��)��v���[`@���K�i^ے�$�	u�i�Oc槢'�	�����am��sٌ0�rƲag;d�j2C�9�X�/o����9��Ⱥ� tՀN�;Qm0�ו�Y�>K��*�	V��0_�tx�)\r�mͣ&�+���]���(���N�ӟ���n�\�ߌ�_�L!½\8��˞+�
l�2�0ߛ�	Ϟ��t�~�5c��%Ҍ�*I�	��N��vqv�`�Y�&Ƨ3
M/�B��I!A0���
L�1�?�X�F�I~�|*esU�S��!-/-��Ί㿀@�H��]a�D���^P�=��^����R5�Oí���_����J���HM$K��v�yQ���0٨���PE����sY}�\��3�Ϲ�+d+Mp�x#��o5�d����V�*�ۋ��Z�V�_b�h�>ʐ��U�;���f_d��zU/�W p�rE8P�3���