BZh91AY&SY	�� _�Px��w߰����P^tF`QD$��=54M�Dm4 �4�F�P�`&F F&&	�bi���B���@z@4�� �@�&d`bba0�!�&�	
z&�I�M5=I��~��M�=4��O�I@���B I�{H>L	����k����xL��V.���V���8`�5���k��l�x�:&I��vDgܾ�$�d���'��\?L�;Jc�,����J�� �=^�l��;F4��.�\�l��b���ɔс_v��p�a;j���9�b��V�1iފ��Պ�%�@�� HgN�o�ne��<�ID���%5S)JM�,�!Є���E&��GIƘ��H`kL�t������J���1�Z5���#���$�G���?�&&j��S�SM���j/šh��w�S(J�^s}���E)�6|7��к4i�m,C1b�g��(��U��q�M�DJV��y�6*r��R^������8�i�⌈#��\�����f�q��P�q�� �[@��2aB^���'�����%×~k>�G-*�k��N��5#�$p�h[�S;��N�65���.I��`�B�ϼh
�68`���:�1dINyS�\�)D(
yf@L�t�����%���y�ZF���t(����!��i�$.8.��0�:a`�v�lP,�8���&!�Bv@�nS9��h$dL2��	�RY�;&�f�pQ�ȃ�a �����7��=��@V�~�aRT	���([���۬��@�(.ը)�{1�D0�$���A���'O/9�.^��̾J�򁙒���!y���H�
A6��