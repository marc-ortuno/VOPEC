BZh91AY&SY�!Z� ߀Px��߰����P~tF`PRS��T�I��Q�j��PG��@昙2h�`��` ���OQT44 �  �9�&L�0�&&��!�0# � �	�AD�ʙ h��zM=K�'�$�A@F�$��$�m%�2�<&�<�
��U���`U�-�^&�Y�7%��6�Agg���}���.����UE*2� �c=gљ2�w
�K4IT������ߑC�Ƙ�U�\a�&����C�T�3����C_M��ԓ,UPj��L�9AL\�YZU�\��z�o�B�	��Ά�o;+��EQmq1*���M��V��
�M�Ta9�D�N5F��.����,d�K.����a���Ɓ��S*��8�r�$��g�f���>UP�B�{�:HNn��)x��ƬV�x��f!�xؠ=��'��!H.�B���=��f�.g�~���1�ا��P���i��sq9ͤDJV��8�ۛ�2���=$ټ��p�WE�,�\K����j�?a��,�0��"aB^ވ���SF�"K���:,�;s�a�Q��״��H�7��`Y��o�Ad:5K¦��
�H�!�h�a�i�TV�C�Z�#	�P5<e��B�0��D$���H��T��P�+�N��7��{2����uĘz0�>�4�e�f^k�|�&��É�z�iڑؘ�����H�ν�P�VZl�ui$�w޿��Ve�vdn7i�%@�+-�B΢"#]��x�E���G��CI �,P��:��\00��l>s�G�D�׼m"l@"�	���)�
��