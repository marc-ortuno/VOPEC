BZh91AY&SY���] �߀Px���߰����Px<���+ABP�SʛSz���4=@OQ� � �5=       		�4�M46�  544d���`F�b0L�`�!4��4=Sjjf#HyM z��&�i���B�$�H@3��E�5f�bF��h�~l�\�I1�0�������q�.���d!2d!2��-҇��:W{L��߼=7�u�"e���NѪuP��F�VT�D庬[���{���ج(3Q<`����5(�Mb��;�kj���R#c=�՚�J- CL��c�ı���6y`UnMʦ�m�X��_�9�L�P�f���ɪ��J�#�%r"h�u�P"����R�$.�	$��
(S0� �=&�AV��Pq*�B�B4��`���0��v@�3LGr
�`��,TY�
��
;�JjLՠCĮk4SVú�tG���%'	�C ���ƨnƣ}��co���lB.}�5���c|>%0U�X��䱕��0�<�M�5�Ξ*1�9ED� Ƒ�p���p� ū.�C�xk������Iٯ-�es�s��%w��֤Ǔ�J�z,4���5b0 g-.����LZ�E��_�	]"��&p����J��2*e@��<�M���x��*������@v�!�ų`��ap�*
���g�|�_���A��ˀ蓠����/�*Z�V�Kϩ�ӗ5�%!/|f��zM�k
��D��_�Jx����D$*ghh��;�L�E]�\+1���(^0(טrȳ��je�}aC�A��3��U�A�P�o�_���F�����iOz۽I=�Nv��PY����hH��X�a�u�nf&�щ��f�>��V���@M4`l`%�}�R�@ѱ�:��l[hLw�������HX�jY2��YJ`Ѕ$�L��l$�0e,�� �t[�H�!hWY���L%/j��;N��F��B|7#0��	�x�5���30if;�b%�Z�p�{Ĝ2��"�͂#:�6���9f^��h�H9&4���qP���7�oP��E��X�@!t�$;�2�?>��7�t�� +��Jb�R�L�V�@2��=� $ͅMW�j+W��u* ���Of�>�:�������$�S	�FC���TO¤|�u�)c0��~�T��ܑN$:7�W@