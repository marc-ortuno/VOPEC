BZh91AY&SYd�� c߀Px��g߰����P�wm���Hez�4Q� �� �  %	��~����@    ����4�L�hh�   s	�L �L&�  L�hH��&��!&�&�!�#�bc����X�$�2�m%�C!��|��`�ƑS;P�����ND���I�܆��$��Rtm�DJ2���F/�_���r�Hk�k(ł�R�ȕŸ%LjN"%**�$Z����P�!�1�j�b��E�T��^���ד��"��I��
a�T4�]�Y;`��.�Y��)���'�g;	5�E6T�ӽ�l�N��<5�� B�C2t��V�vX�O%(�n��LAD�L��"�K�N��q�&Ch0����'Cg�i���5��������O�W�����x��y#��a����!�@�������V��
� �娼Hi[��Ő|N�� ��$���a��c�B��k<8V�(]<Q�vb��s�$TE�Iò����uD��eI`kc�)�(dD�vy�&�+�5�i�qFD���F�32���	������/&%��G�vܘ1����ӷ]=��䍸T�[4>\3��Ԏ�F���
��_a��+/lz��U`ꪚ$�XfhFa���LZ�=��Ea�2�1e$���PjwKm�(�@�S�� �d�c�?�L YVU<L�\�QTt�
a�ZD=f�HZ�.|d�y�9+ݙ�m�`Zf�� ^�3��pjU�!ؑ�1��eIHeS4Ꚅk����eh����Bam/[�pI)��*`��F�!r��"S@���ihZ2y@�f,AMຢ�a�H-��>�P{���b2B,͞�{[[�1wXq��0T+?�w$S�	�O��