BZh91AY&SY��-� �ߔPx��o߰����   Prqg3F�%L&��DS#@zA�h�M4T�&��L�d   � 2d�2@  hi�4d���`F�b0L�`� �i�5S���M'�M����(����H�IP@X�D������,
4��������xLB�ib�jmY�h�s��j���(�ʅ��G�5�*���}̬
ah�n0s�/\���VV����L�>�^ifRH�+!�s>�}p�(T�1�+�=
�B.>��=���9HeXHo�Ή>
v� )`@b+��C�_���x#�t�@Y�"L �YU�U,&j�$)�P�@x���"��J,$�Z�N����Pf�a'[�Nf�66�m��W(G�<��w��$9zPIf�HA�!ݐ "��� ��Cl/R$�6Y�X@UI�[�ٙ�qÔ�)��>��g���i��a�
.4FB���N�'�j��/�8�
�4�{�L,$|�b�^m@�m������?��� �!�@v+�O��P��%)��ω�5�� $k�l-X!�CFp�F�K���KX`�����s8��N�nP�%�]��&�׼`���+⌆�lˑ��^P��� �r�>��ZA�Xcq�iDH*L���ي`�#"!��f�%YL(���V�(�(�tS�o�Mw 9����/�%p�Zf�&B���zD��z7!�	��`Xm(ő �s��2�J$(
y� 	&N:C��`y��O��u�E�Xv�B�G?-�{�h�̜��P�[4au����R8��"�M;��&��٠�	�m�$)2��{#���F��6��	(o?=�n{�E��ߕ0�*�%m� ����A�4���Y`S1�ƥëA4V"���P�1	*{Sܪ�e)^���PT		��)��]��BC;䶔