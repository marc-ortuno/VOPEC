BZh91AY&SY �� }_�Px��߰����P8�s&��X$��?S�${M$ѐ4��2���`RD �    	L��@��<�L��� !�昙2h�`��` ���RH&Hm&�L#҆O$h��zL�N,+�I$&(FBI^��g�B��yKT�x_V=��*F4�����L����kĲ�Ie���T�Xd1p��Ě��cg�{�r)�b��������HSSR4�J��:&�̊JT4��oH�m?��آ��)�1�-E[���M.��Z\�k=�q��u�J���:�;�}.Nz<�5Υw����!2�0�����ߪˁ&b�L`��Hȫ-!�š�ә�L�ԙ I'wGj؅z$h�8yl�T�����dBL�,���HN
{f|Yn�U�!��t У2�e�u�HLPm=������áB���&�x+4�٨�hb�����$�	l�I�#t���p�B�=�CIF�i�5�B�p�w��<���x7^�q���'F�wMX�9/�mHBBKBI P 1�����pps���4x�o2�ĩ�Ȏ�#�,��ȊR ��!B GR*X����:3-*! ��:�o2��>�/�0ɧ/�΄�G]�m���.�'1q�!状��WNkt-D 0��w-F-����+@u\��,Yɳ����Ǫki]ͻR�^A�.�-:����<����9}����,�I~׎0��C�x��M��n�6;Z�_aǼ�-ũKN��ǲB�� ��p��evCQ�^�>�C[T>@U�7����9
ߗ)�6���������(�-�ӂ������d8���@C�Xج����db�C�sn�>Z�uO��5c�����T�n��)I���i��f�mNf�.8귁Ei�=%�@2[��0&LB�^�x��I~�|�esU�S���庻zkc` o��K�Ts��U�����	��7z����P�����2����)S��xD\�5`���Z:��0�f�tl\ZYZ���l]j�ۜ0a|���rl2p��F������8��m`t�Q��rlłQ�ľ�XM�����S�L�l��L�̾ȧϞ�q���5O�.�p� �14