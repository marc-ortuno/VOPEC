BZh91AY&SY�2 @߀Px��o߰����P^sl��V�	$�=��5G�h�4 � s �	������`���`%2!D4�M42  � s �	������`���`$�#B��ɩ<Б����� D��!_	$�"]	�E�W��Y�PƤ�@��y<q��QU#*O���eS%Ÿ����qC61�c��p���cw�p�C��Ɲq8�ܑ�R��&R�D����5�W��ĕ���R6G!x�p
��7a!ɖ�g��}�AJ��<���f[��j�+pvflY��aG���2�=7a�|�5�P,��kV,��L٪e�Mj��d��ZH����#S�+�U[ck\�,)E]�;�9�U���F��t��5v1q�F5�x�Xf%��Y�]g�q.qyVC[m�r�dgYۃl����9˵�[|GY!		-�$�@�����(�MGuw��*�J�� �O�b�F&DAJ
 Њ��jn����6�� % %�W����_���d�2�R��;z���J=EĂ$9I����|��SE��1{�J�o�+��E�4wV�I�� � �Z�,w�N����LZG9�)iʞ��3�ODN`���׃I�/m�ǡ�Ⱥ����9�	�|xiD�־W�v�����i�r|���1H�S�PW$�e��^���SN,�ù�v��*�\e���~	��N�nm�+�1��~��(�[r���uv��::X;w�(��Åz�qko�<:���i�_~n ��}R�O~隲���J3p���S�);�/��v*��lht�I���w1ۇv��",B�Ca�+5�t��ߊ�8�e-�L�:�-1-˟R+�� �0N['˩���
�kN�N.*/��Z���1��%�Y�씩�ψ7D���w_,�������"q�a 98m"-��tp�P��H·�bG���Nw-=KZ�᭬֥��s�=��&&��P5�	�� ˈ}�rE7���53/����Rcd�&AL'�rE8P��2